module collide_top( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [15:0] io_Link_A_X1_In, // @[:@6.4]
  input  [15:0] io_Link_A_X0_In, // @[:@6.4]
  input  [15:0] io_Link_A_Y1_In, // @[:@6.4]
  input  [15:0] io_Link_A_Y0_In, // @[:@6.4]
  input  [15:0] io_Link_A_Z1_In, // @[:@6.4]
  input  [15:0] io_Link_A_Z0_In, // @[:@6.4]
  input  [15:0] io_Link_B_X1_In, // @[:@6.4]
  input  [15:0] io_Link_B_X0_In, // @[:@6.4]
  input  [15:0] io_Link_B_Y1_In, // @[:@6.4]
  input  [15:0] io_Link_B_Y0_In, // @[:@6.4]
  input  [15:0] io_Link_B_Z1_In, // @[:@6.4]
  input  [15:0] io_Link_B_Z0_In, // @[:@6.4]
  output [17:0] io_distance, // @[:@6.4]
  input  [7:0]  io_state // @[:@6.4]
);
  wire [8:0] _T_45; // @[collide_top.scala 49:37:@20.4]
  wire [8:0] Link_A_X1; // @[collide_top.scala 49:44:@21.4]
  wire [8:0] _T_47; // @[collide_top.scala 50:37:@23.4]
  wire [8:0] Link_A_X0; // @[collide_top.scala 50:44:@24.4]
  wire [8:0] _T_49; // @[collide_top.scala 51:37:@26.4]
  wire [8:0] Link_A_Y1; // @[collide_top.scala 51:44:@27.4]
  wire [8:0] _T_51; // @[collide_top.scala 52:37:@29.4]
  wire [8:0] Link_A_Y0; // @[collide_top.scala 52:44:@30.4]
  wire [8:0] _T_53; // @[collide_top.scala 53:37:@32.4]
  wire [8:0] Link_A_Z1; // @[collide_top.scala 53:44:@33.4]
  wire [8:0] _T_55; // @[collide_top.scala 54:37:@35.4]
  wire [8:0] Link_A_Z0; // @[collide_top.scala 54:44:@36.4]
  wire [8:0] _T_57; // @[collide_top.scala 55:37:@38.4]
  wire [8:0] Link_B_X1; // @[collide_top.scala 55:44:@39.4]
  wire [8:0] _T_59; // @[collide_top.scala 56:37:@41.4]
  wire [8:0] Link_B_X0; // @[collide_top.scala 56:44:@42.4]
  wire [8:0] _T_61; // @[collide_top.scala 57:37:@44.4]
  wire [8:0] Link_B_Y1; // @[collide_top.scala 57:44:@45.4]
  wire [8:0] _T_63; // @[collide_top.scala 58:37:@47.4]
  wire [8:0] Link_B_Y0; // @[collide_top.scala 58:44:@48.4]
  wire [8:0] _T_65; // @[collide_top.scala 59:37:@50.4]
  wire [8:0] Link_B_Z1; // @[collide_top.scala 59:44:@51.4]
  wire [8:0] _T_67; // @[collide_top.scala 60:37:@53.4]
  wire [8:0] Link_B_Z0; // @[collide_top.scala 60:44:@54.4]
  reg [8:0] ux; // @[collide_top.scala 64:21:@56.4]
  reg [31:0] _RAND_0;
  reg [8:0] uy; // @[collide_top.scala 65:21:@57.4]
  reg [31:0] _RAND_1;
  reg [8:0] uz; // @[collide_top.scala 66:21:@58.4]
  reg [31:0] _RAND_2;
  reg [8:0] vx; // @[collide_top.scala 67:21:@59.4]
  reg [31:0] _RAND_3;
  reg [8:0] vy; // @[collide_top.scala 68:21:@60.4]
  reg [31:0] _RAND_4;
  reg [8:0] vz; // @[collide_top.scala 69:21:@61.4]
  reg [31:0] _RAND_5;
  reg [8:0] wx; // @[collide_top.scala 70:21:@62.4]
  reg [31:0] _RAND_6;
  reg [8:0] wy; // @[collide_top.scala 71:21:@63.4]
  reg [31:0] _RAND_7;
  reg [8:0] wz; // @[collide_top.scala 72:21:@64.4]
  reg [31:0] _RAND_8;
  reg [17:0] uxux; // @[collide_top.scala 74:23:@65.4]
  reg [31:0] _RAND_9;
  reg [17:0] uyuy; // @[collide_top.scala 75:23:@66.4]
  reg [31:0] _RAND_10;
  reg [17:0] uzuz; // @[collide_top.scala 76:23:@67.4]
  reg [31:0] _RAND_11;
  reg [17:0] uxvx; // @[collide_top.scala 78:23:@68.4]
  reg [31:0] _RAND_12;
  reg [17:0] uyvy; // @[collide_top.scala 79:23:@69.4]
  reg [31:0] _RAND_13;
  reg [17:0] uzvz; // @[collide_top.scala 80:23:@70.4]
  reg [31:0] _RAND_14;
  reg [17:0] vxvx; // @[collide_top.scala 82:23:@71.4]
  reg [31:0] _RAND_15;
  reg [17:0] vyvy; // @[collide_top.scala 83:23:@72.4]
  reg [31:0] _RAND_16;
  reg [17:0] vzvz; // @[collide_top.scala 84:23:@73.4]
  reg [31:0] _RAND_17;
  reg [17:0] uxwx; // @[collide_top.scala 86:23:@74.4]
  reg [31:0] _RAND_18;
  reg [17:0] uywy; // @[collide_top.scala 87:23:@75.4]
  reg [31:0] _RAND_19;
  reg [17:0] uzwz; // @[collide_top.scala 88:23:@76.4]
  reg [31:0] _RAND_20;
  reg [17:0] vxwx; // @[collide_top.scala 90:23:@77.4]
  reg [31:0] _RAND_21;
  reg [17:0] vywy; // @[collide_top.scala 91:23:@78.4]
  reg [31:0] _RAND_22;
  reg [17:0] vzwz; // @[collide_top.scala 92:23:@79.4]
  reg [31:0] _RAND_23;
  reg [17:0] a; // @[collide_top.scala 94:20:@80.4]
  reg [31:0] _RAND_24;
  reg [17:0] b; // @[collide_top.scala 95:20:@81.4]
  reg [31:0] _RAND_25;
  reg [17:0] c; // @[collide_top.scala 96:20:@82.4]
  reg [31:0] _RAND_26;
  reg [17:0] d; // @[collide_top.scala 97:20:@83.4]
  reg [31:0] _RAND_27;
  reg [17:0] e; // @[collide_top.scala 98:20:@84.4]
  reg [31:0] _RAND_28;
  reg [35:0] a_ex; // @[collide_top.scala 100:23:@85.4]
  reg [63:0] _RAND_29;
  reg [35:0] b_ex; // @[collide_top.scala 101:23:@86.4]
  reg [63:0] _RAND_30;
  reg [35:0] c_ex; // @[collide_top.scala 102:23:@87.4]
  reg [63:0] _RAND_31;
  reg [35:0] d_ex; // @[collide_top.scala 103:23:@88.4]
  reg [63:0] _RAND_32;
  reg [35:0] e_ex; // @[collide_top.scala 104:23:@89.4]
  reg [63:0] _RAND_33;
  reg [35:0] ac; // @[collide_top.scala 106:21:@90.4]
  reg [63:0] _RAND_34;
  reg [35:0] bb; // @[collide_top.scala 107:21:@91.4]
  reg [63:0] _RAND_35;
  reg [35:0] be; // @[collide_top.scala 108:21:@92.4]
  reg [63:0] _RAND_36;
  reg [35:0] cd; // @[collide_top.scala 109:21:@93.4]
  reg [63:0] _RAND_37;
  reg [35:0] ae; // @[collide_top.scala 110:21:@94.4]
  reg [63:0] _RAND_38;
  reg [35:0] bd; // @[collide_top.scala 111:21:@95.4]
  reg [63:0] _RAND_39;
  reg [35:0] D_SUB_B; // @[collide_top.scala 123:26:@100.4]
  reg [63:0] _RAND_40;
  reg [35:0] sn_temp; // @[collide_top.scala 125:26:@101.4]
  reg [63:0] _RAND_41;
  reg [35:0] sd_temp; // @[collide_top.scala 126:26:@102.4]
  reg [63:0] _RAND_42;
  reg [35:0] tn_temp; // @[collide_top.scala 127:26:@103.4]
  reg [63:0] _RAND_43;
  reg [35:0] td; // @[collide_top.scala 128:21:@104.4]
  reg [63:0] _RAND_44;
  reg [5:0] sc; // @[collide_top.scala 132:21:@105.4]
  reg [31:0] _RAND_45;
  reg [5:0] tc; // @[collide_top.scala 133:21:@106.4]
  reg [31:0] _RAND_46;
  reg [40:0] sn_calData; // @[collide_top.scala 135:29:@107.4]
  reg [63:0] _RAND_47;
  reg [40:0] sd_calData; // @[collide_top.scala 136:29:@108.4]
  reg [63:0] _RAND_48;
  reg [40:0] tn_calData; // @[collide_top.scala 138:29:@109.4]
  reg [63:0] _RAND_49;
  reg [40:0] td_calData; // @[collide_top.scala 139:29:@110.4]
  reg [63:0] _RAND_50;
  reg [14:0] scux; // @[collide_top.scala 141:23:@111.4]
  reg [31:0] _RAND_51;
  reg [14:0] tcvx; // @[collide_top.scala 142:23:@112.4]
  reg [31:0] _RAND_52;
  reg [14:0] scuy; // @[collide_top.scala 143:23:@113.4]
  reg [31:0] _RAND_53;
  reg [14:0] tcvy; // @[collide_top.scala 144:23:@114.4]
  reg [31:0] _RAND_54;
  reg [14:0] scuz; // @[collide_top.scala 145:23:@115.4]
  reg [31:0] _RAND_55;
  reg [14:0] tcvz; // @[collide_top.scala 146:23:@116.4]
  reg [31:0] _RAND_56;
  reg [8:0] dx; // @[collide_top.scala 148:21:@117.4]
  reg [31:0] _RAND_57;
  reg [8:0] dy; // @[collide_top.scala 149:21:@118.4]
  reg [31:0] _RAND_58;
  reg [8:0] dz; // @[collide_top.scala 150:21:@119.4]
  reg [31:0] _RAND_59;
  reg [17:0] dxdx; // @[collide_top.scala 152:23:@120.4]
  reg [31:0] _RAND_60;
  reg [17:0] dydy; // @[collide_top.scala 153:23:@121.4]
  reg [31:0] _RAND_61;
  reg [17:0] dzdz; // @[collide_top.scala 154:23:@122.4]
  reg [31:0] _RAND_62;
  wire [41:0] _GEN_955; // @[collide_top.scala 185:40:@143.4]
  wire [41:0] _T_152; // @[collide_top.scala 185:40:@143.4]
  wire [40:0] sn_calData_move1; // @[collide_top.scala 163:36:@123.4 collide_top.scala 185:26:@144.4]
  wire  SC_CMP_S1; // @[collide_top.scala 180:39:@135.4]
  wire [41:0] _T_156; // @[collide_top.scala 190:83:@151.4]
  wire [41:0] _T_157; // @[collide_top.scala 190:83:@152.4]
  wire [40:0] _T_158; // @[collide_top.scala 190:83:@153.4]
  wire [40:0] SN_CALDATA_COMPRESS; // @[collide_top.scala 190:35:@154.4]
  wire [41:0] _GEN_956; // @[collide_top.scala 186:49:@145.4]
  wire [41:0] _T_153; // @[collide_top.scala 186:49:@145.4]
  wire [40:0] sn_calData_move2; // @[collide_top.scala 164:36:@124.4 collide_top.scala 186:26:@146.4]
  wire  SC_CMP_S2; // @[collide_top.scala 181:39:@137.4]
  wire [41:0] _GEN_957; // @[collide_top.scala 187:40:@147.4]
  wire [41:0] _T_154; // @[collide_top.scala 187:40:@147.4]
  wire [40:0] tn_calData_move1; // @[collide_top.scala 168:36:@127.4 collide_top.scala 187:26:@148.4]
  wire  TC_CMP_S1; // @[collide_top.scala 182:39:@139.4]
  wire [41:0] _T_165; // @[collide_top.scala 192:83:@161.4]
  wire [41:0] _T_166; // @[collide_top.scala 192:83:@162.4]
  wire [40:0] _T_167; // @[collide_top.scala 192:83:@163.4]
  wire [40:0] TN_CALDATA_COMPRESS; // @[collide_top.scala 192:35:@164.4]
  wire [41:0] _GEN_958; // @[collide_top.scala 188:49:@149.4]
  wire [41:0] _T_155; // @[collide_top.scala 188:49:@149.4]
  wire [40:0] tn_calData_move2; // @[collide_top.scala 169:36:@128.4 collide_top.scala 188:26:@150.4]
  wire  TC_CMP_S2; // @[collide_top.scala 183:39:@141.4]
  wire [6:0] _GEN_959; // @[collide_top.scala 191:45:@156.4]
  wire [6:0] _T_160; // @[collide_top.scala 191:45:@156.4]
  wire [6:0] _T_163; // @[collide_top.scala 191:64:@158.4]
  wire [6:0] _T_164; // @[collide_top.scala 191:27:@159.4]
  wire [6:0] _GEN_961; // @[collide_top.scala 193:45:@166.4]
  wire [6:0] _T_169; // @[collide_top.scala 193:45:@166.4]
  wire [6:0] _T_172; // @[collide_top.scala 193:64:@168.4]
  wire [6:0] _T_173; // @[collide_top.scala 193:27:@169.4]
  wire [36:0] _T_213; // @[collide_top.scala 230:25:@213.4]
  wire [35:0] _T_214; // @[collide_top.scala 230:25:@214.4]
  wire [35:0] AC_SUB_BB; // @[collide_top.scala 230:25:@215.4]
  wire  flag_parallel; // @[collide_top.scala 198:37:@173.4]
  wire [36:0] _T_216; // @[collide_top.scala 231:25:@217.4]
  wire [35:0] _T_217; // @[collide_top.scala 231:25:@218.4]
  wire [35:0] BE_SUB_CD; // @[collide_top.scala 231:25:@219.4]
  wire  Foot1OutofSta; // @[collide_top.scala 199:37:@175.4]
  wire [36:0] _T_183; // @[collide_top.scala 205:47:@180.4]
  wire [35:0] _T_184; // @[collide_top.scala 205:47:@181.4]
  wire [35:0] BE_SUB_CD_SSUB_AC_SUB_BB; // @[collide_top.scala 205:47:@182.4]
  wire  _T_186; // @[collide_top.scala 206:51:@184.4]
  wire  Foot1OutofEnd; // @[collide_top.scala 206:56:@185.4]
  wire  Foot2OutofSta; // @[collide_top.scala 211:35:@188.4]
  wire [36:0] _T_195; // @[collide_top.scala 216:35:@193.4]
  wire [35:0] _T_196; // @[collide_top.scala 216:35:@194.4]
  wire [35:0] TN_TEMP_SUB_TD; // @[collide_top.scala 216:35:@195.4]
  wire  _T_198; // @[collide_top.scala 217:42:@197.4]
  wire  Foot2OutofEnd; // @[collide_top.scala 217:47:@198.4]
  wire  _T_202; // @[collide_top.scala 221:24:@201.4]
  wire  D_CMPB_0; // @[collide_top.scala 221:29:@202.4]
  wire [18:0] _T_207; // @[collide_top.scala 226:22:@206.4]
  wire [17:0] _T_208; // @[collide_top.scala 226:22:@207.4]
  wire [17:0] D_ADD_A; // @[collide_top.scala 226:22:@208.4]
  wire  D_CMPS_nA; // @[collide_top.scala 227:31:@210.4]
  wire [36:0] _T_219; // @[collide_top.scala 232:25:@221.4]
  wire [35:0] _T_220; // @[collide_top.scala 232:25:@222.4]
  wire [35:0] AE_SUB_BD; // @[collide_top.scala 232:25:@223.4]
  wire [36:0] _T_222; // @[collide_top.scala 233:26:@225.4]
  wire [35:0] _T_223; // @[collide_top.scala 233:26:@226.4]
  wire [35:0] E_ADD_B; // @[collide_top.scala 233:26:@227.4]
  wire  _T_226; // @[collide_top.scala 237:36:@230.4]
  wire  D_SUB_B_CMPB_0; // @[collide_top.scala 237:41:@231.4]
  wire [36:0] _T_231; // @[collide_top.scala 242:34:@235.4]
  wire [35:0] _T_232; // @[collide_top.scala 242:34:@236.4]
  wire [35:0] D_SUB_B_ADD_A; // @[collide_top.scala 242:34:@237.4]
  wire  D_SUB_B_CMPS_nA; // @[collide_top.scala 243:43:@239.4]
  reg [17:0] distance_Reg; // @[collide_top.scala 245:31:@242.4]
  reg [31:0] _RAND_63;
  wire  _T_304; // @[collide_top.scala 331:24:@311.6]
  wire [9:0] _T_305; // @[collide_top.scala 333:33:@313.8]
  wire [8:0] _T_306; // @[collide_top.scala 333:33:@314.8]
  wire [8:0] _T_307; // @[collide_top.scala 333:33:@315.8]
  wire [9:0] _T_308; // @[collide_top.scala 334:33:@317.8]
  wire [8:0] _T_309; // @[collide_top.scala 334:33:@318.8]
  wire [8:0] _T_310; // @[collide_top.scala 334:33:@319.8]
  wire [9:0] _T_311; // @[collide_top.scala 335:33:@321.8]
  wire [8:0] _T_312; // @[collide_top.scala 335:33:@322.8]
  wire [8:0] _T_313; // @[collide_top.scala 335:33:@323.8]
  wire [9:0] _T_314; // @[collide_top.scala 337:33:@325.8]
  wire [8:0] _T_315; // @[collide_top.scala 337:33:@326.8]
  wire [8:0] _T_316; // @[collide_top.scala 337:33:@327.8]
  wire [9:0] _T_317; // @[collide_top.scala 338:33:@329.8]
  wire [8:0] _T_318; // @[collide_top.scala 338:33:@330.8]
  wire [8:0] _T_319; // @[collide_top.scala 338:33:@331.8]
  wire [9:0] _T_320; // @[collide_top.scala 339:33:@333.8]
  wire [8:0] _T_321; // @[collide_top.scala 339:33:@334.8]
  wire [8:0] _T_322; // @[collide_top.scala 339:33:@335.8]
  wire [9:0] _T_323; // @[collide_top.scala 341:33:@337.8]
  wire [8:0] _T_324; // @[collide_top.scala 341:33:@338.8]
  wire [8:0] _T_325; // @[collide_top.scala 341:33:@339.8]
  wire [9:0] _T_326; // @[collide_top.scala 342:33:@341.8]
  wire [8:0] _T_327; // @[collide_top.scala 342:33:@342.8]
  wire [8:0] _T_328; // @[collide_top.scala 342:33:@343.8]
  wire [9:0] _T_329; // @[collide_top.scala 343:33:@345.8]
  wire [8:0] _T_330; // @[collide_top.scala 343:33:@346.8]
  wire [8:0] _T_331; // @[collide_top.scala 343:33:@347.8]
  wire  _T_333; // @[collide_top.scala 345:29:@351.8]
  wire [17:0] _T_334; // @[collide_top.scala 347:28:@353.10]
  wire [17:0] _T_335; // @[collide_top.scala 348:28:@355.10]
  wire [17:0] _T_336; // @[collide_top.scala 349:28:@357.10]
  wire [17:0] _T_337; // @[collide_top.scala 350:28:@359.10]
  wire [17:0] _T_338; // @[collide_top.scala 351:28:@361.10]
  wire [17:0] _T_339; // @[collide_top.scala 352:28:@363.10]
  wire [17:0] _T_340; // @[collide_top.scala 353:28:@365.10]
  wire [17:0] _T_341; // @[collide_top.scala 354:28:@367.10]
  wire [17:0] _T_342; // @[collide_top.scala 355:28:@369.10]
  wire [17:0] _T_343; // @[collide_top.scala 356:28:@371.10]
  wire [17:0] _T_344; // @[collide_top.scala 357:28:@373.10]
  wire [17:0] _T_345; // @[collide_top.scala 358:28:@375.10]
  wire [17:0] _T_346; // @[collide_top.scala 359:28:@377.10]
  wire [17:0] _T_347; // @[collide_top.scala 360:28:@379.10]
  wire [17:0] _T_348; // @[collide_top.scala 361:28:@381.10]
  wire  _T_350; // @[collide_top.scala 363:29:@385.10]
  wire [18:0] _T_351; // @[collide_top.scala 365:27:@387.12]
  wire [17:0] _T_352; // @[collide_top.scala 365:27:@388.12]
  wire [17:0] _T_353; // @[collide_top.scala 365:27:@389.12]
  wire [18:0] _T_354; // @[collide_top.scala 365:34:@390.12]
  wire [17:0] _T_355; // @[collide_top.scala 365:34:@391.12]
  wire [17:0] _T_356; // @[collide_top.scala 365:34:@392.12]
  wire [18:0] _T_357; // @[collide_top.scala 366:27:@394.12]
  wire [17:0] _T_358; // @[collide_top.scala 366:27:@395.12]
  wire [17:0] _T_359; // @[collide_top.scala 366:27:@396.12]
  wire [18:0] _T_360; // @[collide_top.scala 366:34:@397.12]
  wire [17:0] _T_361; // @[collide_top.scala 366:34:@398.12]
  wire [17:0] _T_362; // @[collide_top.scala 366:34:@399.12]
  wire [18:0] _T_363; // @[collide_top.scala 367:27:@401.12]
  wire [17:0] _T_364; // @[collide_top.scala 367:27:@402.12]
  wire [17:0] _T_365; // @[collide_top.scala 367:27:@403.12]
  wire [18:0] _T_366; // @[collide_top.scala 367:34:@404.12]
  wire [17:0] _T_367; // @[collide_top.scala 367:34:@405.12]
  wire [17:0] _T_368; // @[collide_top.scala 367:34:@406.12]
  wire [18:0] _T_369; // @[collide_top.scala 368:27:@408.12]
  wire [17:0] _T_370; // @[collide_top.scala 368:27:@409.12]
  wire [17:0] _T_371; // @[collide_top.scala 368:27:@410.12]
  wire [18:0] _T_372; // @[collide_top.scala 368:34:@411.12]
  wire [17:0] _T_373; // @[collide_top.scala 368:34:@412.12]
  wire [17:0] _T_374; // @[collide_top.scala 368:34:@413.12]
  wire [18:0] _T_375; // @[collide_top.scala 369:27:@415.12]
  wire [17:0] _T_376; // @[collide_top.scala 369:27:@416.12]
  wire [17:0] _T_377; // @[collide_top.scala 369:27:@417.12]
  wire [18:0] _T_378; // @[collide_top.scala 369:34:@418.12]
  wire [17:0] _T_379; // @[collide_top.scala 369:34:@419.12]
  wire [17:0] _T_380; // @[collide_top.scala 369:34:@420.12]
  wire  _T_382; // @[collide_top.scala 372:29:@424.12]
  wire [35:0] _T_383; // @[collide_top.scala 374:25:@426.14]
  wire [35:0] _T_384; // @[collide_top.scala 375:25:@428.14]
  wire [35:0] _T_385; // @[collide_top.scala 376:25:@430.14]
  wire [35:0] _T_386; // @[collide_top.scala 377:25:@432.14]
  wire [35:0] _T_387; // @[collide_top.scala 378:25:@434.14]
  wire [35:0] _T_388; // @[collide_top.scala 379:25:@436.14]
  wire  _T_389; // @[collide_top.scala 381:39:@438.14]
  wire [17:0] _T_393; // @[Bitwise.scala 72:12:@440.14]
  wire [17:0] _T_394; // @[collide_top.scala 381:48:@441.14]
  wire [35:0] _T_395; // @[Cat.scala 30:58:@442.14]
  wire [35:0] _T_396; // @[collide_top.scala 381:57:@443.14]
  wire  _T_397; // @[collide_top.scala 382:39:@445.14]
  wire [17:0] _T_401; // @[Bitwise.scala 72:12:@447.14]
  wire [17:0] _T_402; // @[collide_top.scala 382:48:@448.14]
  wire [35:0] _T_403; // @[Cat.scala 30:58:@449.14]
  wire [35:0] _T_404; // @[collide_top.scala 382:57:@450.14]
  wire  _T_405; // @[collide_top.scala 383:39:@452.14]
  wire [17:0] _T_409; // @[Bitwise.scala 72:12:@454.14]
  wire [17:0] _T_410; // @[collide_top.scala 383:48:@455.14]
  wire [35:0] _T_411; // @[Cat.scala 30:58:@456.14]
  wire [35:0] _T_412; // @[collide_top.scala 383:57:@457.14]
  wire [17:0] _T_417; // @[Bitwise.scala 72:12:@461.14]
  wire [17:0] _T_418; // @[collide_top.scala 384:48:@462.14]
  wire [35:0] _T_419; // @[Cat.scala 30:58:@463.14]
  wire [35:0] _T_420; // @[collide_top.scala 384:57:@464.14]
  wire  _T_421; // @[collide_top.scala 385:39:@466.14]
  wire [17:0] _T_425; // @[Bitwise.scala 72:12:@468.14]
  wire [17:0] _T_426; // @[collide_top.scala 385:48:@469.14]
  wire [35:0] _T_427; // @[Cat.scala 30:58:@470.14]
  wire [35:0] _T_428; // @[collide_top.scala 385:57:@471.14]
  wire  _T_430; // @[collide_top.scala 387:29:@475.14]
  wire [36:0] _T_431; // @[collide_top.scala 389:33:@477.16]
  wire [35:0] _T_432; // @[collide_top.scala 389:33:@478.16]
  wire [35:0] _T_433; // @[collide_top.scala 389:33:@479.16]
  wire [36:0] _T_437; // @[collide_top.scala 393:87:@481.16]
  wire [35:0] _T_438; // @[collide_top.scala 393:87:@482.16]
  wire [35:0] _T_439; // @[collide_top.scala 393:87:@483.16]
  wire [35:0] _T_440; // @[collide_top.scala 393:60:@484.16]
  wire [35:0] _T_441; // @[collide_top.scala 392:52:@485.16]
  wire [35:0] _T_442; // @[collide_top.scala 391:31:@486.16]
  wire [35:0] _T_444; // @[collide_top.scala 398:31:@488.16]
  wire [35:0] _T_445; // @[collide_top.scala 403:60:@490.16]
  wire [35:0] _T_446; // @[collide_top.scala 402:52:@491.16]
  wire [35:0] _T_447; // @[collide_top.scala 401:31:@492.16]
  wire [35:0] _T_448; // @[collide_top.scala 410:52:@494.16]
  wire [35:0] _T_449; // @[collide_top.scala 409:44:@495.16]
  wire [35:0] _T_450; // @[collide_top.scala 408:28:@496.16]
  wire  _T_452; // @[collide_top.scala 415:29:@500.16]
  wire [36:0] _T_456; // @[collide_top.scala 420:112:@502.18]
  wire [35:0] _T_457; // @[collide_top.scala 420:112:@503.18]
  wire [35:0] _T_458; // @[collide_top.scala 420:112:@504.18]
  wire [35:0] _T_459; // @[collide_top.scala 420:119:@505.18]
  wire [35:0] _T_460; // @[collide_top.scala 420:92:@506.18]
  wire [35:0] _T_461; // @[collide_top.scala 419:84:@507.18]
  wire [36:0] _T_465; // @[collide_top.scala 424:158:@508.18]
  wire [35:0] _T_466; // @[collide_top.scala 424:158:@509.18]
  wire [35:0] _T_467; // @[collide_top.scala 424:158:@510.18]
  wire [35:0] _T_468; // @[collide_top.scala 424:168:@511.18]
  wire [35:0] _T_469; // @[collide_top.scala 424:132:@512.18]
  wire [35:0] _T_470; // @[collide_top.scala 423:116:@513.18]
  wire [35:0] _T_471; // @[collide_top.scala 426:130:@514.18]
  wire [35:0] _T_472; // @[collide_top.scala 422:84:@515.18]
  wire [35:0] _T_473; // @[collide_top.scala 418:34:@516.18]
  wire [35:0] _T_474; // @[collide_top.scala 431:106:@518.18]
  wire [35:0] _T_476; // @[collide_top.scala 432:143:@519.18]
  wire [35:0] _T_477; // @[collide_top.scala 432:116:@520.18]
  wire [35:0] _T_478; // @[collide_top.scala 431:84:@521.18]
  wire [35:0] _T_482; // @[collide_top.scala 436:124:@524.18]
  wire [35:0] _T_483; // @[collide_top.scala 435:116:@525.18]
  wire [35:0] _T_485; // @[collide_top.scala 434:84:@527.18]
  wire [35:0] _T_486; // @[collide_top.scala 430:34:@528.18]
  wire [36:0] _T_489; // @[collide_top.scala 445:81:@530.18]
  wire [35:0] _T_490; // @[collide_top.scala 445:81:@531.18]
  wire [35:0] _T_491; // @[collide_top.scala 445:81:@532.18]
  wire [35:0] _T_492; // @[collide_top.scala 445:88:@533.18]
  wire [35:0] _T_493; // @[collide_top.scala 445:106:@534.18]
  wire [35:0] _T_494; // @[collide_top.scala 445:60:@535.18]
  wire [35:0] _T_495; // @[collide_top.scala 444:34:@536.18]
  wire [35:0] _T_496; // @[collide_top.scala 448:36:@538.18]
  wire  _T_500; // @[collide_top.scala 454:29:@544.18]
  wire [41:0] _T_501; // @[collide_top.scala 456:82:@546.20]
  wire [41:0] _T_502; // @[collide_top.scala 456:82:@547.20]
  wire [40:0] _T_503; // @[collide_top.scala 456:82:@548.20]
  wire [40:0] _T_504; // @[collide_top.scala 456:34:@549.20]
  wire [5:0] SC_COMPRESS; // @[collide_top.scala 165:31:@125.4 collide_top.scala 191:21:@160.4]
  wire [6:0] _GEN_963; // @[collide_top.scala 457:50:@551.20]
  wire [6:0] _T_505; // @[collide_top.scala 457:50:@551.20]
  wire [7:0] _T_508; // @[collide_top.scala 457:77:@553.20]
  wire [6:0] _T_509; // @[collide_top.scala 457:77:@554.20]
  wire [6:0] _T_510; // @[collide_top.scala 457:26:@555.20]
  wire [41:0] _T_511; // @[collide_top.scala 459:82:@557.20]
  wire [41:0] _T_512; // @[collide_top.scala 459:82:@558.20]
  wire [40:0] _T_513; // @[collide_top.scala 459:82:@559.20]
  wire [40:0] _T_514; // @[collide_top.scala 459:34:@560.20]
  wire [5:0] TC_COMPRESS; // @[collide_top.scala 170:31:@129.4 collide_top.scala 193:21:@170.4]
  wire [6:0] _GEN_965; // @[collide_top.scala 460:50:@562.20]
  wire [6:0] _T_515; // @[collide_top.scala 460:50:@562.20]
  wire [7:0] _T_518; // @[collide_top.scala 460:77:@564.20]
  wire [6:0] _T_519; // @[collide_top.scala 460:77:@565.20]
  wire [6:0] _T_520; // @[collide_top.scala 460:26:@566.20]
  wire  _T_522; // @[collide_top.scala 463:29:@570.20]
  wire  _T_544; // @[collide_top.scala 471:29:@596.22]
  wire  _T_566; // @[collide_top.scala 479:29:@622.24]
  wire [6:0] _T_567; // @[collide_top.scala 481:28:@624.26]
  wire [8:0] _GEN_975; // @[collide_top.scala 481:28:@625.26]
  wire [15:0] _T_568; // @[collide_top.scala 481:28:@625.26]
  wire [14:0] _T_569; // @[collide_top.scala 481:28:@626.26]
  wire [14:0] _T_570; // @[collide_top.scala 481:28:@627.26]
  wire [6:0] _T_571; // @[collide_top.scala 482:28:@629.26]
  wire [8:0] _GEN_976; // @[collide_top.scala 482:28:@630.26]
  wire [15:0] _T_572; // @[collide_top.scala 482:28:@630.26]
  wire [14:0] _T_573; // @[collide_top.scala 482:28:@631.26]
  wire [14:0] _T_574; // @[collide_top.scala 482:28:@632.26]
  wire [15:0] _T_576; // @[collide_top.scala 483:28:@635.26]
  wire [14:0] _T_577; // @[collide_top.scala 483:28:@636.26]
  wire [14:0] _T_578; // @[collide_top.scala 483:28:@637.26]
  wire [15:0] _T_580; // @[collide_top.scala 484:28:@640.26]
  wire [14:0] _T_581; // @[collide_top.scala 484:28:@641.26]
  wire [14:0] _T_582; // @[collide_top.scala 484:28:@642.26]
  wire [15:0] _T_584; // @[collide_top.scala 485:28:@645.26]
  wire [14:0] _T_585; // @[collide_top.scala 485:28:@646.26]
  wire [14:0] _T_586; // @[collide_top.scala 485:28:@647.26]
  wire [15:0] _T_588; // @[collide_top.scala 486:28:@650.26]
  wire [14:0] _T_589; // @[collide_top.scala 486:28:@651.26]
  wire [14:0] _T_590; // @[collide_top.scala 486:28:@652.26]
  wire  _T_592; // @[collide_top.scala 488:29:@656.26]
  wire [8:0] _T_593; // @[collide_top.scala 490:32:@658.28]
  wire [8:0] _T_594; // @[collide_top.scala 490:39:@659.28]
  wire [9:0] _T_595; // @[collide_top.scala 490:26:@660.28]
  wire [8:0] _T_596; // @[collide_top.scala 490:26:@661.28]
  wire [8:0] _T_597; // @[collide_top.scala 490:26:@662.28]
  wire [8:0] _T_598; // @[collide_top.scala 490:52:@663.28]
  wire [8:0] _T_599; // @[collide_top.scala 490:59:@664.28]
  wire [9:0] _T_600; // @[collide_top.scala 490:46:@665.28]
  wire [8:0] _T_601; // @[collide_top.scala 490:46:@666.28]
  wire [8:0] _T_602; // @[collide_top.scala 490:46:@667.28]
  wire [8:0] _T_603; // @[collide_top.scala 491:32:@669.28]
  wire [8:0] _T_604; // @[collide_top.scala 491:39:@670.28]
  wire [9:0] _T_605; // @[collide_top.scala 491:26:@671.28]
  wire [8:0] _T_606; // @[collide_top.scala 491:26:@672.28]
  wire [8:0] _T_607; // @[collide_top.scala 491:26:@673.28]
  wire [8:0] _T_608; // @[collide_top.scala 491:52:@674.28]
  wire [8:0] _T_609; // @[collide_top.scala 491:59:@675.28]
  wire [9:0] _T_610; // @[collide_top.scala 491:46:@676.28]
  wire [8:0] _T_611; // @[collide_top.scala 491:46:@677.28]
  wire [8:0] _T_612; // @[collide_top.scala 491:46:@678.28]
  wire [8:0] _T_613; // @[collide_top.scala 492:32:@680.28]
  wire [8:0] _T_614; // @[collide_top.scala 492:39:@681.28]
  wire [9:0] _T_615; // @[collide_top.scala 492:26:@682.28]
  wire [8:0] _T_616; // @[collide_top.scala 492:26:@683.28]
  wire [8:0] _T_617; // @[collide_top.scala 492:26:@684.28]
  wire [8:0] _T_618; // @[collide_top.scala 492:52:@685.28]
  wire [8:0] _T_619; // @[collide_top.scala 492:59:@686.28]
  wire [9:0] _T_620; // @[collide_top.scala 492:46:@687.28]
  wire [8:0] _T_621; // @[collide_top.scala 492:46:@688.28]
  wire [8:0] _T_622; // @[collide_top.scala 492:46:@689.28]
  wire  _T_624; // @[collide_top.scala 494:29:@693.28]
  wire [17:0] _T_625; // @[collide_top.scala 496:28:@695.30]
  wire [17:0] _T_626; // @[collide_top.scala 497:28:@697.30]
  wire [17:0] _T_627; // @[collide_top.scala 498:28:@699.30]
  wire  _T_629; // @[collide_top.scala 500:29:@703.30]
  wire [18:0] _T_630; // @[collide_top.scala 502:38:@705.32]
  wire [17:0] _T_631; // @[collide_top.scala 502:38:@706.32]
  wire [17:0] _T_632; // @[collide_top.scala 502:38:@707.32]
  wire [18:0] _T_633; // @[collide_top.scala 502:45:@708.32]
  wire [17:0] _T_634; // @[collide_top.scala 502:45:@709.32]
  wire [17:0] _T_635; // @[collide_top.scala 502:45:@710.32]
  wire  _T_637; // @[collide_top.scala 504:29:@714.32]
  wire [17:0] _GEN_0; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_1; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_2; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_3; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_4; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_5; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_6; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_7; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_8; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_9; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_10; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_11; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_12; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_13; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_14; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_15; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_16; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_17; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_18; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_19; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_20; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_21; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_22; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_23; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_24; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_25; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_26; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_27; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_28; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_29; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_30; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_31; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_32; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_33; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_34; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_35; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_36; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_37; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_38; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_39; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_40; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_41; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_42; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_43; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_44; // @[collide_top.scala 505:9:@715.32]
  wire [35:0] _GEN_45; // @[collide_top.scala 505:9:@715.32]
  wire [5:0] _GEN_46; // @[collide_top.scala 505:9:@715.32]
  wire [5:0] _GEN_47; // @[collide_top.scala 505:9:@715.32]
  wire [40:0] _GEN_48; // @[collide_top.scala 505:9:@715.32]
  wire [40:0] _GEN_49; // @[collide_top.scala 505:9:@715.32]
  wire [40:0] _GEN_50; // @[collide_top.scala 505:9:@715.32]
  wire [14:0] _GEN_51; // @[collide_top.scala 505:9:@715.32]
  wire [14:0] _GEN_52; // @[collide_top.scala 505:9:@715.32]
  wire [14:0] _GEN_53; // @[collide_top.scala 505:9:@715.32]
  wire [14:0] _GEN_54; // @[collide_top.scala 505:9:@715.32]
  wire [14:0] _GEN_55; // @[collide_top.scala 505:9:@715.32]
  wire [14:0] _GEN_56; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_57; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_58; // @[collide_top.scala 505:9:@715.32]
  wire [8:0] _GEN_59; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_60; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_61; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_62; // @[collide_top.scala 505:9:@715.32]
  wire [17:0] _GEN_63; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_64; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_65; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_66; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_67; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_68; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_69; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_70; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_71; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_72; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_73; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_74; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_75; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_76; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_77; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_78; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_79; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_80; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_81; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_82; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_83; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_84; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_85; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_86; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_87; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_88; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_89; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_90; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_91; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_92; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_93; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_94; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_95; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_96; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_97; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_98; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_99; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_100; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_101; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_102; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_103; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_104; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_105; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_106; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_107; // @[collide_top.scala 501:9:@704.30]
  wire [35:0] _GEN_108; // @[collide_top.scala 501:9:@704.30]
  wire [5:0] _GEN_109; // @[collide_top.scala 501:9:@704.30]
  wire [5:0] _GEN_110; // @[collide_top.scala 501:9:@704.30]
  wire [40:0] _GEN_111; // @[collide_top.scala 501:9:@704.30]
  wire [40:0] _GEN_112; // @[collide_top.scala 501:9:@704.30]
  wire [40:0] _GEN_113; // @[collide_top.scala 501:9:@704.30]
  wire [14:0] _GEN_114; // @[collide_top.scala 501:9:@704.30]
  wire [14:0] _GEN_115; // @[collide_top.scala 501:9:@704.30]
  wire [14:0] _GEN_116; // @[collide_top.scala 501:9:@704.30]
  wire [14:0] _GEN_117; // @[collide_top.scala 501:9:@704.30]
  wire [14:0] _GEN_118; // @[collide_top.scala 501:9:@704.30]
  wire [14:0] _GEN_119; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_120; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_121; // @[collide_top.scala 501:9:@704.30]
  wire [8:0] _GEN_122; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_123; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_124; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_125; // @[collide_top.scala 501:9:@704.30]
  wire [17:0] _GEN_126; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_127; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_128; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_129; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_130; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_131; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_132; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_133; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_134; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_135; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_136; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_137; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_138; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_139; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_140; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_141; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_142; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_143; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_144; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_145; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_146; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_147; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_148; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_149; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_150; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_151; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_152; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_153; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_154; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_155; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_156; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_157; // @[collide_top.scala 495:9:@694.28]
  wire [17:0] _GEN_158; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_159; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_160; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_161; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_162; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_163; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_164; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_165; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_166; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_167; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_168; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_169; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_170; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_171; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_172; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_173; // @[collide_top.scala 495:9:@694.28]
  wire [35:0] _GEN_174; // @[collide_top.scala 495:9:@694.28]
  wire [5:0] _GEN_175; // @[collide_top.scala 495:9:@694.28]
  wire [5:0] _GEN_176; // @[collide_top.scala 495:9:@694.28]
  wire [40:0] _GEN_177; // @[collide_top.scala 495:9:@694.28]
  wire [40:0] _GEN_178; // @[collide_top.scala 495:9:@694.28]
  wire [40:0] _GEN_179; // @[collide_top.scala 495:9:@694.28]
  wire [14:0] _GEN_180; // @[collide_top.scala 495:9:@694.28]
  wire [14:0] _GEN_181; // @[collide_top.scala 495:9:@694.28]
  wire [14:0] _GEN_182; // @[collide_top.scala 495:9:@694.28]
  wire [14:0] _GEN_183; // @[collide_top.scala 495:9:@694.28]
  wire [14:0] _GEN_184; // @[collide_top.scala 495:9:@694.28]
  wire [14:0] _GEN_185; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_186; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_187; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_188; // @[collide_top.scala 495:9:@694.28]
  wire [8:0] _GEN_189; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_190; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_191; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_192; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_193; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_194; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_195; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_196; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_197; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_198; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_199; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_200; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_201; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_202; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_203; // @[collide_top.scala 489:9:@657.26]
  wire [8:0] _GEN_204; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_205; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_206; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_207; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_208; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_209; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_210; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_211; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_212; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_213; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_214; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_215; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_216; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_217; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_218; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_219; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_220; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_221; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_222; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_223; // @[collide_top.scala 489:9:@657.26]
  wire [17:0] _GEN_224; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_225; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_226; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_227; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_228; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_229; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_230; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_231; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_232; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_233; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_234; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_235; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_236; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_237; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_238; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_239; // @[collide_top.scala 489:9:@657.26]
  wire [35:0] _GEN_240; // @[collide_top.scala 489:9:@657.26]
  wire [5:0] _GEN_241; // @[collide_top.scala 489:9:@657.26]
  wire [5:0] _GEN_242; // @[collide_top.scala 489:9:@657.26]
  wire [40:0] _GEN_243; // @[collide_top.scala 489:9:@657.26]
  wire [40:0] _GEN_244; // @[collide_top.scala 489:9:@657.26]
  wire [40:0] _GEN_245; // @[collide_top.scala 489:9:@657.26]
  wire [14:0] _GEN_246; // @[collide_top.scala 489:9:@657.26]
  wire [14:0] _GEN_247; // @[collide_top.scala 489:9:@657.26]
  wire [14:0] _GEN_248; // @[collide_top.scala 489:9:@657.26]
  wire [14:0] _GEN_249; // @[collide_top.scala 489:9:@657.26]
  wire [14:0] _GEN_250; // @[collide_top.scala 489:9:@657.26]
  wire [14:0] _GEN_251; // @[collide_top.scala 489:9:@657.26]
  wire [14:0] _GEN_252; // @[collide_top.scala 480:9:@623.24]
  wire [14:0] _GEN_253; // @[collide_top.scala 480:9:@623.24]
  wire [14:0] _GEN_254; // @[collide_top.scala 480:9:@623.24]
  wire [14:0] _GEN_255; // @[collide_top.scala 480:9:@623.24]
  wire [14:0] _GEN_256; // @[collide_top.scala 480:9:@623.24]
  wire [14:0] _GEN_257; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_258; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_259; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_260; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_261; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_262; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_263; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_264; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_265; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_266; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_267; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_268; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_269; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_270; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_271; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_272; // @[collide_top.scala 480:9:@623.24]
  wire [8:0] _GEN_273; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_274; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_275; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_276; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_277; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_278; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_279; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_280; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_281; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_282; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_283; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_284; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_285; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_286; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_287; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_288; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_289; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_290; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_291; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_292; // @[collide_top.scala 480:9:@623.24]
  wire [17:0] _GEN_293; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_294; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_295; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_296; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_297; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_298; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_299; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_300; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_301; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_302; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_303; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_304; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_305; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_306; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_307; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_308; // @[collide_top.scala 480:9:@623.24]
  wire [35:0] _GEN_309; // @[collide_top.scala 480:9:@623.24]
  wire [5:0] _GEN_310; // @[collide_top.scala 480:9:@623.24]
  wire [5:0] _GEN_311; // @[collide_top.scala 480:9:@623.24]
  wire [40:0] _GEN_312; // @[collide_top.scala 480:9:@623.24]
  wire [40:0] _GEN_313; // @[collide_top.scala 480:9:@623.24]
  wire [40:0] _GEN_314; // @[collide_top.scala 480:9:@623.24]
  wire [40:0] _GEN_315; // @[collide_top.scala 472:9:@597.22]
  wire [6:0] _GEN_316; // @[collide_top.scala 472:9:@597.22]
  wire [40:0] _GEN_317; // @[collide_top.scala 472:9:@597.22]
  wire [6:0] _GEN_318; // @[collide_top.scala 472:9:@597.22]
  wire [14:0] _GEN_319; // @[collide_top.scala 472:9:@597.22]
  wire [14:0] _GEN_320; // @[collide_top.scala 472:9:@597.22]
  wire [14:0] _GEN_321; // @[collide_top.scala 472:9:@597.22]
  wire [14:0] _GEN_322; // @[collide_top.scala 472:9:@597.22]
  wire [14:0] _GEN_323; // @[collide_top.scala 472:9:@597.22]
  wire [14:0] _GEN_324; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_325; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_326; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_327; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_328; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_329; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_330; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_331; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_332; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_333; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_334; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_335; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_336; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_337; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_338; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_339; // @[collide_top.scala 472:9:@597.22]
  wire [8:0] _GEN_340; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_341; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_342; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_343; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_344; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_345; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_346; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_347; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_348; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_349; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_350; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_351; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_352; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_353; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_354; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_355; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_356; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_357; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_358; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_359; // @[collide_top.scala 472:9:@597.22]
  wire [17:0] _GEN_360; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_361; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_362; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_363; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_364; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_365; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_366; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_367; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_368; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_369; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_370; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_371; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_372; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_373; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_374; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_375; // @[collide_top.scala 472:9:@597.22]
  wire [35:0] _GEN_376; // @[collide_top.scala 472:9:@597.22]
  wire [40:0] _GEN_377; // @[collide_top.scala 472:9:@597.22]
  wire [40:0] _GEN_378; // @[collide_top.scala 472:9:@597.22]
  wire [40:0] _GEN_379; // @[collide_top.scala 464:9:@571.20]
  wire [6:0] _GEN_380; // @[collide_top.scala 464:9:@571.20]
  wire [40:0] _GEN_381; // @[collide_top.scala 464:9:@571.20]
  wire [6:0] _GEN_382; // @[collide_top.scala 464:9:@571.20]
  wire [14:0] _GEN_383; // @[collide_top.scala 464:9:@571.20]
  wire [14:0] _GEN_384; // @[collide_top.scala 464:9:@571.20]
  wire [14:0] _GEN_385; // @[collide_top.scala 464:9:@571.20]
  wire [14:0] _GEN_386; // @[collide_top.scala 464:9:@571.20]
  wire [14:0] _GEN_387; // @[collide_top.scala 464:9:@571.20]
  wire [14:0] _GEN_388; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_389; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_390; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_391; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_392; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_393; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_394; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_395; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_396; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_397; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_398; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_399; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_400; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_401; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_402; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_403; // @[collide_top.scala 464:9:@571.20]
  wire [8:0] _GEN_404; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_405; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_406; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_407; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_408; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_409; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_410; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_411; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_412; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_413; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_414; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_415; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_416; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_417; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_418; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_419; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_420; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_421; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_422; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_423; // @[collide_top.scala 464:9:@571.20]
  wire [17:0] _GEN_424; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_425; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_426; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_427; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_428; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_429; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_430; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_431; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_432; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_433; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_434; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_435; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_436; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_437; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_438; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_439; // @[collide_top.scala 464:9:@571.20]
  wire [35:0] _GEN_440; // @[collide_top.scala 464:9:@571.20]
  wire [40:0] _GEN_441; // @[collide_top.scala 464:9:@571.20]
  wire [40:0] _GEN_442; // @[collide_top.scala 464:9:@571.20]
  wire [40:0] _GEN_443; // @[collide_top.scala 455:9:@545.18]
  wire [6:0] _GEN_444; // @[collide_top.scala 455:9:@545.18]
  wire [40:0] _GEN_445; // @[collide_top.scala 455:9:@545.18]
  wire [6:0] _GEN_446; // @[collide_top.scala 455:9:@545.18]
  wire [14:0] _GEN_447; // @[collide_top.scala 455:9:@545.18]
  wire [14:0] _GEN_448; // @[collide_top.scala 455:9:@545.18]
  wire [14:0] _GEN_449; // @[collide_top.scala 455:9:@545.18]
  wire [14:0] _GEN_450; // @[collide_top.scala 455:9:@545.18]
  wire [14:0] _GEN_451; // @[collide_top.scala 455:9:@545.18]
  wire [14:0] _GEN_452; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_453; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_454; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_455; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_456; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_457; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_458; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_459; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_460; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_461; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_462; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_463; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_464; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_465; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_466; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_467; // @[collide_top.scala 455:9:@545.18]
  wire [8:0] _GEN_468; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_469; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_470; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_471; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_472; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_473; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_474; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_475; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_476; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_477; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_478; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_479; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_480; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_481; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_482; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_483; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_484; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_485; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_486; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_487; // @[collide_top.scala 455:9:@545.18]
  wire [17:0] _GEN_488; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_489; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_490; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_491; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_492; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_493; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_494; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_495; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_496; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_497; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_498; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_499; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_500; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_501; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_502; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_503; // @[collide_top.scala 455:9:@545.18]
  wire [35:0] _GEN_504; // @[collide_top.scala 455:9:@545.18]
  wire [40:0] _GEN_505; // @[collide_top.scala 455:9:@545.18]
  wire [40:0] _GEN_506; // @[collide_top.scala 455:9:@545.18]
  wire [40:0] _GEN_507; // @[collide_top.scala 416:9:@501.16]
  wire [40:0] _GEN_508; // @[collide_top.scala 416:9:@501.16]
  wire [40:0] _GEN_509; // @[collide_top.scala 416:9:@501.16]
  wire [40:0] _GEN_510; // @[collide_top.scala 416:9:@501.16]
  wire [6:0] _GEN_511; // @[collide_top.scala 416:9:@501.16]
  wire [6:0] _GEN_512; // @[collide_top.scala 416:9:@501.16]
  wire [14:0] _GEN_513; // @[collide_top.scala 416:9:@501.16]
  wire [14:0] _GEN_514; // @[collide_top.scala 416:9:@501.16]
  wire [14:0] _GEN_515; // @[collide_top.scala 416:9:@501.16]
  wire [14:0] _GEN_516; // @[collide_top.scala 416:9:@501.16]
  wire [14:0] _GEN_517; // @[collide_top.scala 416:9:@501.16]
  wire [14:0] _GEN_518; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_519; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_520; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_521; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_522; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_523; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_524; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_525; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_526; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_527; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_528; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_529; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_530; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_531; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_532; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_533; // @[collide_top.scala 416:9:@501.16]
  wire [8:0] _GEN_534; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_535; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_536; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_537; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_538; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_539; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_540; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_541; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_542; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_543; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_544; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_545; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_546; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_547; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_548; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_549; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_550; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_551; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_552; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_553; // @[collide_top.scala 416:9:@501.16]
  wire [17:0] _GEN_554; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_555; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_556; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_557; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_558; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_559; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_560; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_561; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_562; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_563; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_564; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_565; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_566; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_567; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_568; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_569; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_570; // @[collide_top.scala 416:9:@501.16]
  wire [35:0] _GEN_571; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_572; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_573; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_574; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_575; // @[collide_top.scala 388:9:@476.14]
  wire [40:0] _GEN_576; // @[collide_top.scala 388:9:@476.14]
  wire [40:0] _GEN_577; // @[collide_top.scala 388:9:@476.14]
  wire [40:0] _GEN_578; // @[collide_top.scala 388:9:@476.14]
  wire [40:0] _GEN_579; // @[collide_top.scala 388:9:@476.14]
  wire [6:0] _GEN_580; // @[collide_top.scala 388:9:@476.14]
  wire [6:0] _GEN_581; // @[collide_top.scala 388:9:@476.14]
  wire [14:0] _GEN_582; // @[collide_top.scala 388:9:@476.14]
  wire [14:0] _GEN_583; // @[collide_top.scala 388:9:@476.14]
  wire [14:0] _GEN_584; // @[collide_top.scala 388:9:@476.14]
  wire [14:0] _GEN_585; // @[collide_top.scala 388:9:@476.14]
  wire [14:0] _GEN_586; // @[collide_top.scala 388:9:@476.14]
  wire [14:0] _GEN_587; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_588; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_589; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_590; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_591; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_592; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_593; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_594; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_595; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_596; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_597; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_598; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_599; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_600; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_601; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_602; // @[collide_top.scala 388:9:@476.14]
  wire [8:0] _GEN_603; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_604; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_605; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_606; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_607; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_608; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_609; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_610; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_611; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_612; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_613; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_614; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_615; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_616; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_617; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_618; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_619; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_620; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_621; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_622; // @[collide_top.scala 388:9:@476.14]
  wire [17:0] _GEN_623; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_624; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_625; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_626; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_627; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_628; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_629; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_630; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_631; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_632; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_633; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_634; // @[collide_top.scala 388:9:@476.14]
  wire [35:0] _GEN_635; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_636; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_637; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_638; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_639; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_640; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_641; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_642; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_643; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_644; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_645; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_646; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_647; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_648; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_649; // @[collide_top.scala 373:9:@425.12]
  wire [35:0] _GEN_650; // @[collide_top.scala 373:9:@425.12]
  wire [40:0] _GEN_651; // @[collide_top.scala 373:9:@425.12]
  wire [40:0] _GEN_652; // @[collide_top.scala 373:9:@425.12]
  wire [40:0] _GEN_653; // @[collide_top.scala 373:9:@425.12]
  wire [40:0] _GEN_654; // @[collide_top.scala 373:9:@425.12]
  wire [6:0] _GEN_655; // @[collide_top.scala 373:9:@425.12]
  wire [6:0] _GEN_656; // @[collide_top.scala 373:9:@425.12]
  wire [14:0] _GEN_657; // @[collide_top.scala 373:9:@425.12]
  wire [14:0] _GEN_658; // @[collide_top.scala 373:9:@425.12]
  wire [14:0] _GEN_659; // @[collide_top.scala 373:9:@425.12]
  wire [14:0] _GEN_660; // @[collide_top.scala 373:9:@425.12]
  wire [14:0] _GEN_661; // @[collide_top.scala 373:9:@425.12]
  wire [14:0] _GEN_662; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_663; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_664; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_665; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_666; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_667; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_668; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_669; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_670; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_671; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_672; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_673; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_674; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_675; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_676; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_677; // @[collide_top.scala 373:9:@425.12]
  wire [8:0] _GEN_678; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_679; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_680; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_681; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_682; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_683; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_684; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_685; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_686; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_687; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_688; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_689; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_690; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_691; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_692; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_693; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_694; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_695; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_696; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_697; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_698; // @[collide_top.scala 373:9:@425.12]
  wire [17:0] _GEN_699; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_700; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_701; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_702; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_703; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_704; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_705; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_706; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_707; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_708; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_709; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_710; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_711; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_712; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_713; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_714; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_715; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_716; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_717; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_718; // @[collide_top.scala 364:9:@386.10]
  wire [35:0] _GEN_719; // @[collide_top.scala 364:9:@386.10]
  wire [40:0] _GEN_720; // @[collide_top.scala 364:9:@386.10]
  wire [40:0] _GEN_721; // @[collide_top.scala 364:9:@386.10]
  wire [40:0] _GEN_722; // @[collide_top.scala 364:9:@386.10]
  wire [40:0] _GEN_723; // @[collide_top.scala 364:9:@386.10]
  wire [6:0] _GEN_724; // @[collide_top.scala 364:9:@386.10]
  wire [6:0] _GEN_725; // @[collide_top.scala 364:9:@386.10]
  wire [14:0] _GEN_726; // @[collide_top.scala 364:9:@386.10]
  wire [14:0] _GEN_727; // @[collide_top.scala 364:9:@386.10]
  wire [14:0] _GEN_728; // @[collide_top.scala 364:9:@386.10]
  wire [14:0] _GEN_729; // @[collide_top.scala 364:9:@386.10]
  wire [14:0] _GEN_730; // @[collide_top.scala 364:9:@386.10]
  wire [14:0] _GEN_731; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_732; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_733; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_734; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_735; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_736; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_737; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_738; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_739; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_740; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_741; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_742; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_743; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_744; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_745; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_746; // @[collide_top.scala 364:9:@386.10]
  wire [8:0] _GEN_747; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_748; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_749; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_750; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_751; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_752; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_753; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_754; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_755; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_756; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_757; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_758; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_759; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_760; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_761; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_762; // @[collide_top.scala 364:9:@386.10]
  wire [17:0] _GEN_763; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_764; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_765; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_766; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_767; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_768; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_769; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_770; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_771; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_772; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_773; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_774; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_775; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_776; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_777; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_778; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_779; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_780; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_781; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_782; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_783; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_784; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_785; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_786; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_787; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_788; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_789; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_790; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_791; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_792; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_793; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_794; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_795; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_796; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_797; // @[collide_top.scala 346:9:@352.8]
  wire [35:0] _GEN_798; // @[collide_top.scala 346:9:@352.8]
  wire [40:0] _GEN_799; // @[collide_top.scala 346:9:@352.8]
  wire [40:0] _GEN_800; // @[collide_top.scala 346:9:@352.8]
  wire [40:0] _GEN_801; // @[collide_top.scala 346:9:@352.8]
  wire [40:0] _GEN_802; // @[collide_top.scala 346:9:@352.8]
  wire [6:0] _GEN_803; // @[collide_top.scala 346:9:@352.8]
  wire [6:0] _GEN_804; // @[collide_top.scala 346:9:@352.8]
  wire [14:0] _GEN_805; // @[collide_top.scala 346:9:@352.8]
  wire [14:0] _GEN_806; // @[collide_top.scala 346:9:@352.8]
  wire [14:0] _GEN_807; // @[collide_top.scala 346:9:@352.8]
  wire [14:0] _GEN_808; // @[collide_top.scala 346:9:@352.8]
  wire [14:0] _GEN_809; // @[collide_top.scala 346:9:@352.8]
  wire [14:0] _GEN_810; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_811; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_812; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_813; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_814; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_815; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_816; // @[collide_top.scala 346:9:@352.8]
  wire [17:0] _GEN_817; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_818; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_819; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_820; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_821; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_822; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_823; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_824; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_825; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_826; // @[collide_top.scala 346:9:@352.8]
  wire [8:0] _GEN_827; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_828; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_829; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_830; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_831; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_832; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_833; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_834; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_835; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_836; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_837; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_838; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_839; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_840; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_841; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_842; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_843; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_844; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_845; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_846; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_847; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_848; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_849; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_850; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_851; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_852; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_853; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_854; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_855; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_856; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_857; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_858; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_859; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_860; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_861; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_862; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_863; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_864; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_865; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_866; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_867; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_868; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_869; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_870; // @[collide_top.scala 332:9:@312.6]
  wire [35:0] _GEN_871; // @[collide_top.scala 332:9:@312.6]
  wire [40:0] _GEN_872; // @[collide_top.scala 332:9:@312.6]
  wire [40:0] _GEN_873; // @[collide_top.scala 332:9:@312.6]
  wire [40:0] _GEN_874; // @[collide_top.scala 332:9:@312.6]
  wire [40:0] _GEN_875; // @[collide_top.scala 332:9:@312.6]
  wire [6:0] _GEN_876; // @[collide_top.scala 332:9:@312.6]
  wire [6:0] _GEN_877; // @[collide_top.scala 332:9:@312.6]
  wire [14:0] _GEN_878; // @[collide_top.scala 332:9:@312.6]
  wire [14:0] _GEN_879; // @[collide_top.scala 332:9:@312.6]
  wire [14:0] _GEN_880; // @[collide_top.scala 332:9:@312.6]
  wire [14:0] _GEN_881; // @[collide_top.scala 332:9:@312.6]
  wire [14:0] _GEN_882; // @[collide_top.scala 332:9:@312.6]
  wire [14:0] _GEN_883; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_884; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_885; // @[collide_top.scala 332:9:@312.6]
  wire [8:0] _GEN_886; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_887; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_888; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_889; // @[collide_top.scala 332:9:@312.6]
  wire [17:0] _GEN_890; // @[collide_top.scala 332:9:@312.6]
  wire [6:0] _GEN_936; // @[collide_top.scala 250:1:@244.4]
  wire [6:0] _GEN_937; // @[collide_top.scala 250:1:@244.4]
  assign _T_45 = io_Link_A_X1_In[13:5]; // @[collide_top.scala 49:37:@20.4]
  assign Link_A_X1 = $signed(_T_45); // @[collide_top.scala 49:44:@21.4]
  assign _T_47 = io_Link_A_X0_In[13:5]; // @[collide_top.scala 50:37:@23.4]
  assign Link_A_X0 = $signed(_T_47); // @[collide_top.scala 50:44:@24.4]
  assign _T_49 = io_Link_A_Y1_In[13:5]; // @[collide_top.scala 51:37:@26.4]
  assign Link_A_Y1 = $signed(_T_49); // @[collide_top.scala 51:44:@27.4]
  assign _T_51 = io_Link_A_Y0_In[13:5]; // @[collide_top.scala 52:37:@29.4]
  assign Link_A_Y0 = $signed(_T_51); // @[collide_top.scala 52:44:@30.4]
  assign _T_53 = io_Link_A_Z1_In[13:5]; // @[collide_top.scala 53:37:@32.4]
  assign Link_A_Z1 = $signed(_T_53); // @[collide_top.scala 53:44:@33.4]
  assign _T_55 = io_Link_A_Z0_In[13:5]; // @[collide_top.scala 54:37:@35.4]
  assign Link_A_Z0 = $signed(_T_55); // @[collide_top.scala 54:44:@36.4]
  assign _T_57 = io_Link_B_X1_In[13:5]; // @[collide_top.scala 55:37:@38.4]
  assign Link_B_X1 = $signed(_T_57); // @[collide_top.scala 55:44:@39.4]
  assign _T_59 = io_Link_B_X0_In[13:5]; // @[collide_top.scala 56:37:@41.4]
  assign Link_B_X0 = $signed(_T_59); // @[collide_top.scala 56:44:@42.4]
  assign _T_61 = io_Link_B_Y1_In[13:5]; // @[collide_top.scala 57:37:@44.4]
  assign Link_B_Y1 = $signed(_T_61); // @[collide_top.scala 57:44:@45.4]
  assign _T_63 = io_Link_B_Y0_In[13:5]; // @[collide_top.scala 58:37:@47.4]
  assign Link_B_Y0 = $signed(_T_63); // @[collide_top.scala 58:44:@48.4]
  assign _T_65 = io_Link_B_Z1_In[13:5]; // @[collide_top.scala 59:37:@50.4]
  assign Link_B_Z1 = $signed(_T_65); // @[collide_top.scala 59:44:@51.4]
  assign _T_67 = io_Link_B_Z0_In[13:5]; // @[collide_top.scala 60:37:@53.4]
  assign Link_B_Z0 = $signed(_T_67); // @[collide_top.scala 60:44:@54.4]
  assign _GEN_955 = {{1'd0}, sn_calData}; // @[collide_top.scala 185:40:@143.4]
  assign _T_152 = _GEN_955 << 1; // @[collide_top.scala 185:40:@143.4]
  assign sn_calData_move1 = _T_152[40:0]; // @[collide_top.scala 163:36:@123.4 collide_top.scala 185:26:@144.4]
  assign SC_CMP_S1 = sn_calData_move1 < sd_calData; // @[collide_top.scala 180:39:@135.4]
  assign _T_156 = sn_calData_move1 - sd_calData; // @[collide_top.scala 190:83:@151.4]
  assign _T_157 = $unsigned(_T_156); // @[collide_top.scala 190:83:@152.4]
  assign _T_158 = _T_157[40:0]; // @[collide_top.scala 190:83:@153.4]
  assign SN_CALDATA_COMPRESS = SC_CMP_S1 ? sn_calData_move1 : _T_158; // @[collide_top.scala 190:35:@154.4]
  assign _GEN_956 = {{1'd0}, SN_CALDATA_COMPRESS}; // @[collide_top.scala 186:49:@145.4]
  assign _T_153 = _GEN_956 << 1; // @[collide_top.scala 186:49:@145.4]
  assign sn_calData_move2 = _T_153[40:0]; // @[collide_top.scala 164:36:@124.4 collide_top.scala 186:26:@146.4]
  assign SC_CMP_S2 = sn_calData_move2 < sd_calData; // @[collide_top.scala 181:39:@137.4]
  assign _GEN_957 = {{1'd0}, tn_calData}; // @[collide_top.scala 187:40:@147.4]
  assign _T_154 = _GEN_957 << 1; // @[collide_top.scala 187:40:@147.4]
  assign tn_calData_move1 = _T_154[40:0]; // @[collide_top.scala 168:36:@127.4 collide_top.scala 187:26:@148.4]
  assign TC_CMP_S1 = tn_calData_move1 < td_calData; // @[collide_top.scala 182:39:@139.4]
  assign _T_165 = tn_calData_move1 - td_calData; // @[collide_top.scala 192:83:@161.4]
  assign _T_166 = $unsigned(_T_165); // @[collide_top.scala 192:83:@162.4]
  assign _T_167 = _T_166[40:0]; // @[collide_top.scala 192:83:@163.4]
  assign TN_CALDATA_COMPRESS = TC_CMP_S1 ? tn_calData_move1 : _T_167; // @[collide_top.scala 192:35:@164.4]
  assign _GEN_958 = {{1'd0}, TN_CALDATA_COMPRESS}; // @[collide_top.scala 188:49:@149.4]
  assign _T_155 = _GEN_958 << 1; // @[collide_top.scala 188:49:@149.4]
  assign tn_calData_move2 = _T_155[40:0]; // @[collide_top.scala 169:36:@128.4 collide_top.scala 188:26:@150.4]
  assign TC_CMP_S2 = tn_calData_move2 < td_calData; // @[collide_top.scala 183:39:@141.4]
  assign _GEN_959 = {{1'd0}, sc}; // @[collide_top.scala 191:45:@156.4]
  assign _T_160 = _GEN_959 << 1; // @[collide_top.scala 191:45:@156.4]
  assign _T_163 = _T_160 | 7'h1; // @[collide_top.scala 191:64:@158.4]
  assign _T_164 = SC_CMP_S1 ? _T_160 : _T_163; // @[collide_top.scala 191:27:@159.4]
  assign _GEN_961 = {{1'd0}, tc}; // @[collide_top.scala 193:45:@166.4]
  assign _T_169 = _GEN_961 << 1; // @[collide_top.scala 193:45:@166.4]
  assign _T_172 = _T_169 | 7'h1; // @[collide_top.scala 193:64:@168.4]
  assign _T_173 = TC_CMP_S1 ? _T_169 : _T_172; // @[collide_top.scala 193:27:@169.4]
  assign _T_213 = $signed(ac) - $signed(bb); // @[collide_top.scala 230:25:@213.4]
  assign _T_214 = $signed(ac) - $signed(bb); // @[collide_top.scala 230:25:@214.4]
  assign AC_SUB_BB = $signed(_T_214); // @[collide_top.scala 230:25:@215.4]
  assign flag_parallel = $signed(AC_SUB_BB) == $signed(36'sh0); // @[collide_top.scala 198:37:@173.4]
  assign _T_216 = $signed(be) - $signed(cd); // @[collide_top.scala 231:25:@217.4]
  assign _T_217 = $signed(be) - $signed(cd); // @[collide_top.scala 231:25:@218.4]
  assign BE_SUB_CD = $signed(_T_217); // @[collide_top.scala 231:25:@219.4]
  assign Foot1OutofSta = BE_SUB_CD[35]; // @[collide_top.scala 199:37:@175.4]
  assign _T_183 = $signed(BE_SUB_CD) - $signed(AC_SUB_BB); // @[collide_top.scala 205:47:@180.4]
  assign _T_184 = $signed(BE_SUB_CD) - $signed(AC_SUB_BB); // @[collide_top.scala 205:47:@181.4]
  assign BE_SUB_CD_SSUB_AC_SUB_BB = $signed(_T_184); // @[collide_top.scala 205:47:@182.4]
  assign _T_186 = BE_SUB_CD_SSUB_AC_SUB_BB[35]; // @[collide_top.scala 206:51:@184.4]
  assign Foot1OutofEnd = _T_186 == 1'h0; // @[collide_top.scala 206:56:@185.4]
  assign Foot2OutofSta = tn_temp[35]; // @[collide_top.scala 211:35:@188.4]
  assign _T_195 = $signed(tn_temp) - $signed(td); // @[collide_top.scala 216:35:@193.4]
  assign _T_196 = $signed(tn_temp) - $signed(td); // @[collide_top.scala 216:35:@194.4]
  assign TN_TEMP_SUB_TD = $signed(_T_196); // @[collide_top.scala 216:35:@195.4]
  assign _T_198 = TN_TEMP_SUB_TD[35]; // @[collide_top.scala 217:42:@197.4]
  assign Foot2OutofEnd = _T_198 == 1'h0; // @[collide_top.scala 217:47:@198.4]
  assign _T_202 = d[17]; // @[collide_top.scala 221:24:@201.4]
  assign D_CMPB_0 = _T_202 == 1'h0; // @[collide_top.scala 221:29:@202.4]
  assign _T_207 = $signed(d) + $signed(a); // @[collide_top.scala 226:22:@206.4]
  assign _T_208 = $signed(d) + $signed(a); // @[collide_top.scala 226:22:@207.4]
  assign D_ADD_A = $signed(_T_208); // @[collide_top.scala 226:22:@208.4]
  assign D_CMPS_nA = D_ADD_A[17]; // @[collide_top.scala 227:31:@210.4]
  assign _T_219 = $signed(ae) - $signed(bd); // @[collide_top.scala 232:25:@221.4]
  assign _T_220 = $signed(ae) - $signed(bd); // @[collide_top.scala 232:25:@222.4]
  assign AE_SUB_BD = $signed(_T_220); // @[collide_top.scala 232:25:@223.4]
  assign _T_222 = $signed(e_ex) + $signed(b_ex); // @[collide_top.scala 233:26:@225.4]
  assign _T_223 = $signed(e_ex) + $signed(b_ex); // @[collide_top.scala 233:26:@226.4]
  assign E_ADD_B = $signed(_T_223); // @[collide_top.scala 233:26:@227.4]
  assign _T_226 = D_SUB_B[35]; // @[collide_top.scala 237:36:@230.4]
  assign D_SUB_B_CMPB_0 = _T_226 == 1'h0; // @[collide_top.scala 237:41:@231.4]
  assign _T_231 = $signed(D_SUB_B) + $signed(a_ex); // @[collide_top.scala 242:34:@235.4]
  assign _T_232 = $signed(D_SUB_B) + $signed(a_ex); // @[collide_top.scala 242:34:@236.4]
  assign D_SUB_B_ADD_A = $signed(_T_232); // @[collide_top.scala 242:34:@237.4]
  assign D_SUB_B_CMPS_nA = D_SUB_B_ADD_A[35]; // @[collide_top.scala 243:43:@239.4]
  assign _T_304 = io_state == 8'hb; // @[collide_top.scala 331:24:@311.6]
  assign _T_305 = $signed(Link_A_X1) - $signed(Link_A_X0); // @[collide_top.scala 333:33:@313.8]
  assign _T_306 = $signed(Link_A_X1) - $signed(Link_A_X0); // @[collide_top.scala 333:33:@314.8]
  assign _T_307 = $signed(_T_306); // @[collide_top.scala 333:33:@315.8]
  assign _T_308 = $signed(Link_A_Y1) - $signed(Link_A_Y0); // @[collide_top.scala 334:33:@317.8]
  assign _T_309 = $signed(Link_A_Y1) - $signed(Link_A_Y0); // @[collide_top.scala 334:33:@318.8]
  assign _T_310 = $signed(_T_309); // @[collide_top.scala 334:33:@319.8]
  assign _T_311 = $signed(Link_A_Z1) - $signed(Link_A_Z0); // @[collide_top.scala 335:33:@321.8]
  assign _T_312 = $signed(Link_A_Z1) - $signed(Link_A_Z0); // @[collide_top.scala 335:33:@322.8]
  assign _T_313 = $signed(_T_312); // @[collide_top.scala 335:33:@323.8]
  assign _T_314 = $signed(Link_B_X1) - $signed(Link_B_X0); // @[collide_top.scala 337:33:@325.8]
  assign _T_315 = $signed(Link_B_X1) - $signed(Link_B_X0); // @[collide_top.scala 337:33:@326.8]
  assign _T_316 = $signed(_T_315); // @[collide_top.scala 337:33:@327.8]
  assign _T_317 = $signed(Link_B_Y1) - $signed(Link_B_Y0); // @[collide_top.scala 338:33:@329.8]
  assign _T_318 = $signed(Link_B_Y1) - $signed(Link_B_Y0); // @[collide_top.scala 338:33:@330.8]
  assign _T_319 = $signed(_T_318); // @[collide_top.scala 338:33:@331.8]
  assign _T_320 = $signed(Link_B_Z1) - $signed(Link_B_Z0); // @[collide_top.scala 339:33:@333.8]
  assign _T_321 = $signed(Link_B_Z1) - $signed(Link_B_Z0); // @[collide_top.scala 339:33:@334.8]
  assign _T_322 = $signed(_T_321); // @[collide_top.scala 339:33:@335.8]
  assign _T_323 = $signed(Link_A_X0) - $signed(Link_B_X0); // @[collide_top.scala 341:33:@337.8]
  assign _T_324 = $signed(Link_A_X0) - $signed(Link_B_X0); // @[collide_top.scala 341:33:@338.8]
  assign _T_325 = $signed(_T_324); // @[collide_top.scala 341:33:@339.8]
  assign _T_326 = $signed(Link_A_Y0) - $signed(Link_B_Y0); // @[collide_top.scala 342:33:@341.8]
  assign _T_327 = $signed(Link_A_Y0) - $signed(Link_B_Y0); // @[collide_top.scala 342:33:@342.8]
  assign _T_328 = $signed(_T_327); // @[collide_top.scala 342:33:@343.8]
  assign _T_329 = $signed(Link_A_Z0) - $signed(Link_B_Z0); // @[collide_top.scala 343:33:@345.8]
  assign _T_330 = $signed(Link_A_Z0) - $signed(Link_B_Z0); // @[collide_top.scala 343:33:@346.8]
  assign _T_331 = $signed(_T_330); // @[collide_top.scala 343:33:@347.8]
  assign _T_333 = io_state == 8'hc; // @[collide_top.scala 345:29:@351.8]
  assign _T_334 = $signed(ux) * $signed(ux); // @[collide_top.scala 347:28:@353.10]
  assign _T_335 = $signed(uy) * $signed(uy); // @[collide_top.scala 348:28:@355.10]
  assign _T_336 = $signed(uz) * $signed(uz); // @[collide_top.scala 349:28:@357.10]
  assign _T_337 = $signed(ux) * $signed(vx); // @[collide_top.scala 350:28:@359.10]
  assign _T_338 = $signed(uy) * $signed(vy); // @[collide_top.scala 351:28:@361.10]
  assign _T_339 = $signed(uz) * $signed(vz); // @[collide_top.scala 352:28:@363.10]
  assign _T_340 = $signed(vx) * $signed(vx); // @[collide_top.scala 353:28:@365.10]
  assign _T_341 = $signed(vy) * $signed(vy); // @[collide_top.scala 354:28:@367.10]
  assign _T_342 = $signed(vz) * $signed(vz); // @[collide_top.scala 355:28:@369.10]
  assign _T_343 = $signed(ux) * $signed(wx); // @[collide_top.scala 356:28:@371.10]
  assign _T_344 = $signed(uy) * $signed(wy); // @[collide_top.scala 357:28:@373.10]
  assign _T_345 = $signed(uz) * $signed(wz); // @[collide_top.scala 358:28:@375.10]
  assign _T_346 = $signed(vx) * $signed(wx); // @[collide_top.scala 359:28:@377.10]
  assign _T_347 = $signed(vy) * $signed(wy); // @[collide_top.scala 360:28:@379.10]
  assign _T_348 = $signed(vz) * $signed(wz); // @[collide_top.scala 361:28:@381.10]
  assign _T_350 = io_state == 8'hd; // @[collide_top.scala 363:29:@385.10]
  assign _T_351 = $signed(uxux) + $signed(uyuy); // @[collide_top.scala 365:27:@387.12]
  assign _T_352 = $signed(uxux) + $signed(uyuy); // @[collide_top.scala 365:27:@388.12]
  assign _T_353 = $signed(_T_352); // @[collide_top.scala 365:27:@389.12]
  assign _T_354 = $signed(_T_353) + $signed(uzuz); // @[collide_top.scala 365:34:@390.12]
  assign _T_355 = $signed(_T_353) + $signed(uzuz); // @[collide_top.scala 365:34:@391.12]
  assign _T_356 = $signed(_T_355); // @[collide_top.scala 365:34:@392.12]
  assign _T_357 = $signed(uxvx) + $signed(uyvy); // @[collide_top.scala 366:27:@394.12]
  assign _T_358 = $signed(uxvx) + $signed(uyvy); // @[collide_top.scala 366:27:@395.12]
  assign _T_359 = $signed(_T_358); // @[collide_top.scala 366:27:@396.12]
  assign _T_360 = $signed(_T_359) + $signed(uzvz); // @[collide_top.scala 366:34:@397.12]
  assign _T_361 = $signed(_T_359) + $signed(uzvz); // @[collide_top.scala 366:34:@398.12]
  assign _T_362 = $signed(_T_361); // @[collide_top.scala 366:34:@399.12]
  assign _T_363 = $signed(vxvx) + $signed(vyvy); // @[collide_top.scala 367:27:@401.12]
  assign _T_364 = $signed(vxvx) + $signed(vyvy); // @[collide_top.scala 367:27:@402.12]
  assign _T_365 = $signed(_T_364); // @[collide_top.scala 367:27:@403.12]
  assign _T_366 = $signed(_T_365) + $signed(vzvz); // @[collide_top.scala 367:34:@404.12]
  assign _T_367 = $signed(_T_365) + $signed(vzvz); // @[collide_top.scala 367:34:@405.12]
  assign _T_368 = $signed(_T_367); // @[collide_top.scala 367:34:@406.12]
  assign _T_369 = $signed(uxwx) + $signed(uywy); // @[collide_top.scala 368:27:@408.12]
  assign _T_370 = $signed(uxwx) + $signed(uywy); // @[collide_top.scala 368:27:@409.12]
  assign _T_371 = $signed(_T_370); // @[collide_top.scala 368:27:@410.12]
  assign _T_372 = $signed(_T_371) + $signed(uzwz); // @[collide_top.scala 368:34:@411.12]
  assign _T_373 = $signed(_T_371) + $signed(uzwz); // @[collide_top.scala 368:34:@412.12]
  assign _T_374 = $signed(_T_373); // @[collide_top.scala 368:34:@413.12]
  assign _T_375 = $signed(vxwx) + $signed(vywy); // @[collide_top.scala 369:27:@415.12]
  assign _T_376 = $signed(vxwx) + $signed(vywy); // @[collide_top.scala 369:27:@416.12]
  assign _T_377 = $signed(_T_376); // @[collide_top.scala 369:27:@417.12]
  assign _T_378 = $signed(_T_377) + $signed(vzwz); // @[collide_top.scala 369:34:@418.12]
  assign _T_379 = $signed(_T_377) + $signed(vzwz); // @[collide_top.scala 369:34:@419.12]
  assign _T_380 = $signed(_T_379); // @[collide_top.scala 369:34:@420.12]
  assign _T_382 = io_state == 8'he; // @[collide_top.scala 372:29:@424.12]
  assign _T_383 = $signed(a) * $signed(c); // @[collide_top.scala 374:25:@426.14]
  assign _T_384 = $signed(b) * $signed(b); // @[collide_top.scala 375:25:@428.14]
  assign _T_385 = $signed(b) * $signed(e); // @[collide_top.scala 376:25:@430.14]
  assign _T_386 = $signed(c) * $signed(d); // @[collide_top.scala 377:25:@432.14]
  assign _T_387 = $signed(a) * $signed(e); // @[collide_top.scala 378:25:@434.14]
  assign _T_388 = $signed(b) * $signed(d); // @[collide_top.scala 379:25:@436.14]
  assign _T_389 = a[17]; // @[collide_top.scala 381:39:@438.14]
  assign _T_393 = _T_389 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12:@440.14]
  assign _T_394 = $unsigned(a); // @[collide_top.scala 381:48:@441.14]
  assign _T_395 = {_T_393,_T_394}; // @[Cat.scala 30:58:@442.14]
  assign _T_396 = $signed(_T_395); // @[collide_top.scala 381:57:@443.14]
  assign _T_397 = b[17]; // @[collide_top.scala 382:39:@445.14]
  assign _T_401 = _T_397 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12:@447.14]
  assign _T_402 = $unsigned(b); // @[collide_top.scala 382:48:@448.14]
  assign _T_403 = {_T_401,_T_402}; // @[Cat.scala 30:58:@449.14]
  assign _T_404 = $signed(_T_403); // @[collide_top.scala 382:57:@450.14]
  assign _T_405 = c[17]; // @[collide_top.scala 383:39:@452.14]
  assign _T_409 = _T_405 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12:@454.14]
  assign _T_410 = $unsigned(c); // @[collide_top.scala 383:48:@455.14]
  assign _T_411 = {_T_409,_T_410}; // @[Cat.scala 30:58:@456.14]
  assign _T_412 = $signed(_T_411); // @[collide_top.scala 383:57:@457.14]
  assign _T_417 = _T_202 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12:@461.14]
  assign _T_418 = $unsigned(d); // @[collide_top.scala 384:48:@462.14]
  assign _T_419 = {_T_417,_T_418}; // @[Cat.scala 30:58:@463.14]
  assign _T_420 = $signed(_T_419); // @[collide_top.scala 384:57:@464.14]
  assign _T_421 = e[17]; // @[collide_top.scala 385:39:@466.14]
  assign _T_425 = _T_421 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12:@468.14]
  assign _T_426 = $unsigned(e); // @[collide_top.scala 385:48:@469.14]
  assign _T_427 = {_T_425,_T_426}; // @[Cat.scala 30:58:@470.14]
  assign _T_428 = $signed(_T_427); // @[collide_top.scala 385:57:@471.14]
  assign _T_430 = io_state == 8'hf; // @[collide_top.scala 387:29:@475.14]
  assign _T_431 = $signed(d_ex) - $signed(b_ex); // @[collide_top.scala 389:33:@477.16]
  assign _T_432 = $signed(d_ex) - $signed(b_ex); // @[collide_top.scala 389:33:@478.16]
  assign _T_433 = $signed(_T_432); // @[collide_top.scala 389:33:@479.16]
  assign _T_437 = $signed(AC_SUB_BB) - $signed(36'sh1); // @[collide_top.scala 393:87:@481.16]
  assign _T_438 = $signed(AC_SUB_BB) - $signed(36'sh1); // @[collide_top.scala 393:87:@482.16]
  assign _T_439 = $signed(_T_438); // @[collide_top.scala 393:87:@483.16]
  assign _T_440 = Foot1OutofEnd ? $signed(_T_439) : $signed(BE_SUB_CD); // @[collide_top.scala 393:60:@484.16]
  assign _T_441 = Foot1OutofSta ? $signed(36'sh0) : $signed(_T_440); // @[collide_top.scala 392:52:@485.16]
  assign _T_442 = flag_parallel ? $signed(36'sh0) : $signed(_T_441); // @[collide_top.scala 391:31:@486.16]
  assign _T_444 = flag_parallel ? $signed(36'sh64) : $signed(AC_SUB_BB); // @[collide_top.scala 398:31:@488.16]
  assign _T_445 = Foot1OutofEnd ? $signed(E_ADD_B) : $signed(AE_SUB_BD); // @[collide_top.scala 403:60:@490.16]
  assign _T_446 = Foot1OutofSta ? $signed(e_ex) : $signed(_T_445); // @[collide_top.scala 402:52:@491.16]
  assign _T_447 = flag_parallel ? $signed(e_ex) : $signed(_T_446); // @[collide_top.scala 401:31:@492.16]
  assign _T_448 = Foot1OutofEnd ? $signed(c_ex) : $signed(AC_SUB_BB); // @[collide_top.scala 410:52:@494.16]
  assign _T_449 = Foot1OutofSta ? $signed(c_ex) : $signed(_T_448); // @[collide_top.scala 409:44:@495.16]
  assign _T_450 = flag_parallel ? $signed(c_ex) : $signed(_T_449); // @[collide_top.scala 408:28:@496.16]
  assign _T_452 = io_state == 8'h10; // @[collide_top.scala 415:29:@500.16]
  assign _T_456 = $signed(36'sh0) - $signed(d_ex); // @[collide_top.scala 420:112:@502.18]
  assign _T_457 = $signed(36'sh0) - $signed(d_ex); // @[collide_top.scala 420:112:@503.18]
  assign _T_458 = $signed(_T_457); // @[collide_top.scala 420:112:@504.18]
  assign _T_459 = $unsigned(_T_458); // @[collide_top.scala 420:119:@505.18]
  assign _T_460 = D_CMPS_nA ? 36'h63 : _T_459; // @[collide_top.scala 420:92:@506.18]
  assign _T_461 = D_CMPB_0 ? 36'h0 : _T_460; // @[collide_top.scala 419:84:@507.18]
  assign _T_465 = $signed(36'sh0) - $signed(D_SUB_B); // @[collide_top.scala 424:158:@508.18]
  assign _T_466 = $signed(36'sh0) - $signed(D_SUB_B); // @[collide_top.scala 424:158:@509.18]
  assign _T_467 = $signed(_T_466); // @[collide_top.scala 424:158:@510.18]
  assign _T_468 = $unsigned(_T_467); // @[collide_top.scala 424:168:@511.18]
  assign _T_469 = D_SUB_B_CMPS_nA ? 36'h63 : _T_468; // @[collide_top.scala 424:132:@512.18]
  assign _T_470 = D_SUB_B_CMPB_0 ? 36'h0 : _T_469; // @[collide_top.scala 423:116:@513.18]
  assign _T_471 = $unsigned(sn_temp); // @[collide_top.scala 426:130:@514.18]
  assign _T_472 = Foot2OutofEnd ? _T_470 : _T_471; // @[collide_top.scala 422:84:@515.18]
  assign _T_473 = Foot2OutofSta ? _T_461 : _T_472; // @[collide_top.scala 418:34:@516.18]
  assign _T_474 = $unsigned(sd_temp); // @[collide_top.scala 431:106:@518.18]
  assign _T_476 = $unsigned(a_ex); // @[collide_top.scala 432:143:@519.18]
  assign _T_477 = D_CMPS_nA ? 36'h64 : _T_476; // @[collide_top.scala 432:116:@520.18]
  assign _T_478 = D_CMPB_0 ? _T_474 : _T_477; // @[collide_top.scala 431:84:@521.18]
  assign _T_482 = D_SUB_B_CMPS_nA ? 36'h64 : _T_476; // @[collide_top.scala 436:124:@524.18]
  assign _T_483 = D_SUB_B_CMPB_0 ? _T_474 : _T_482; // @[collide_top.scala 435:116:@525.18]
  assign _T_485 = Foot2OutofEnd ? _T_483 : _T_474; // @[collide_top.scala 434:84:@527.18]
  assign _T_486 = Foot2OutofSta ? _T_478 : _T_485; // @[collide_top.scala 430:34:@528.18]
  assign _T_489 = $signed(td) - $signed(36'sh1); // @[collide_top.scala 445:81:@530.18]
  assign _T_490 = $signed(td) - $signed(36'sh1); // @[collide_top.scala 445:81:@531.18]
  assign _T_491 = $signed(_T_490); // @[collide_top.scala 445:81:@532.18]
  assign _T_492 = $unsigned(_T_491); // @[collide_top.scala 445:88:@533.18]
  assign _T_493 = $unsigned(tn_temp); // @[collide_top.scala 445:106:@534.18]
  assign _T_494 = Foot2OutofEnd ? _T_492 : _T_493; // @[collide_top.scala 445:60:@535.18]
  assign _T_495 = Foot2OutofSta ? 36'h0 : _T_494; // @[collide_top.scala 444:34:@536.18]
  assign _T_496 = $unsigned(td); // @[collide_top.scala 448:36:@538.18]
  assign _T_500 = io_state == 8'h11; // @[collide_top.scala 454:29:@544.18]
  assign _T_501 = sn_calData_move2 - sd_calData; // @[collide_top.scala 456:82:@546.20]
  assign _T_502 = $unsigned(_T_501); // @[collide_top.scala 456:82:@547.20]
  assign _T_503 = _T_502[40:0]; // @[collide_top.scala 456:82:@548.20]
  assign _T_504 = SC_CMP_S2 ? sn_calData_move2 : _T_503; // @[collide_top.scala 456:34:@549.20]
  assign SC_COMPRESS = _T_164[5:0]; // @[collide_top.scala 165:31:@125.4 collide_top.scala 191:21:@160.4]
  assign _GEN_963 = {{1'd0}, SC_COMPRESS}; // @[collide_top.scala 457:50:@551.20]
  assign _T_505 = _GEN_963 << 1; // @[collide_top.scala 457:50:@551.20]
  assign _T_508 = _T_505 + 7'h1; // @[collide_top.scala 457:77:@553.20]
  assign _T_509 = _T_505 + 7'h1; // @[collide_top.scala 457:77:@554.20]
  assign _T_510 = SC_CMP_S2 ? _T_505 : _T_509; // @[collide_top.scala 457:26:@555.20]
  assign _T_511 = tn_calData_move2 - td_calData; // @[collide_top.scala 459:82:@557.20]
  assign _T_512 = $unsigned(_T_511); // @[collide_top.scala 459:82:@558.20]
  assign _T_513 = _T_512[40:0]; // @[collide_top.scala 459:82:@559.20]
  assign _T_514 = TC_CMP_S2 ? tn_calData_move2 : _T_513; // @[collide_top.scala 459:34:@560.20]
  assign TC_COMPRESS = _T_173[5:0]; // @[collide_top.scala 170:31:@129.4 collide_top.scala 193:21:@170.4]
  assign _GEN_965 = {{1'd0}, TC_COMPRESS}; // @[collide_top.scala 460:50:@562.20]
  assign _T_515 = _GEN_965 << 1; // @[collide_top.scala 460:50:@562.20]
  assign _T_518 = _T_515 + 7'h1; // @[collide_top.scala 460:77:@564.20]
  assign _T_519 = _T_515 + 7'h1; // @[collide_top.scala 460:77:@565.20]
  assign _T_520 = TC_CMP_S2 ? _T_515 : _T_519; // @[collide_top.scala 460:26:@566.20]
  assign _T_522 = io_state == 8'h12; // @[collide_top.scala 463:29:@570.20]
  assign _T_544 = io_state == 8'h13; // @[collide_top.scala 471:29:@596.22]
  assign _T_566 = io_state == 8'h14; // @[collide_top.scala 479:29:@622.24]
  assign _T_567 = {1'b0,$signed(sc)}; // @[collide_top.scala 481:28:@624.26]
  assign _GEN_975 = {{2{_T_567[6]}},_T_567}; // @[collide_top.scala 481:28:@625.26]
  assign _T_568 = $signed(ux) * $signed(_GEN_975); // @[collide_top.scala 481:28:@625.26]
  assign _T_569 = _T_568[14:0]; // @[collide_top.scala 481:28:@626.26]
  assign _T_570 = $signed(_T_569); // @[collide_top.scala 481:28:@627.26]
  assign _T_571 = {1'b0,$signed(tc)}; // @[collide_top.scala 482:28:@629.26]
  assign _GEN_976 = {{2{_T_571[6]}},_T_571}; // @[collide_top.scala 482:28:@630.26]
  assign _T_572 = $signed(vx) * $signed(_GEN_976); // @[collide_top.scala 482:28:@630.26]
  assign _T_573 = _T_572[14:0]; // @[collide_top.scala 482:28:@631.26]
  assign _T_574 = $signed(_T_573); // @[collide_top.scala 482:28:@632.26]
  assign _T_576 = $signed(uy) * $signed(_GEN_975); // @[collide_top.scala 483:28:@635.26]
  assign _T_577 = _T_576[14:0]; // @[collide_top.scala 483:28:@636.26]
  assign _T_578 = $signed(_T_577); // @[collide_top.scala 483:28:@637.26]
  assign _T_580 = $signed(vy) * $signed(_GEN_976); // @[collide_top.scala 484:28:@640.26]
  assign _T_581 = _T_580[14:0]; // @[collide_top.scala 484:28:@641.26]
  assign _T_582 = $signed(_T_581); // @[collide_top.scala 484:28:@642.26]
  assign _T_584 = $signed(uz) * $signed(_GEN_975); // @[collide_top.scala 485:28:@645.26]
  assign _T_585 = _T_584[14:0]; // @[collide_top.scala 485:28:@646.26]
  assign _T_586 = $signed(_T_585); // @[collide_top.scala 485:28:@647.26]
  assign _T_588 = $signed(vz) * $signed(_GEN_976); // @[collide_top.scala 486:28:@650.26]
  assign _T_589 = _T_588[14:0]; // @[collide_top.scala 486:28:@651.26]
  assign _T_590 = $signed(_T_589); // @[collide_top.scala 486:28:@652.26]
  assign _T_592 = io_state == 8'h15; // @[collide_top.scala 488:29:@656.26]
  assign _T_593 = scux[14:6]; // @[collide_top.scala 490:32:@658.28]
  assign _T_594 = $signed(_T_593); // @[collide_top.scala 490:39:@659.28]
  assign _T_595 = $signed(wx) + $signed(_T_594); // @[collide_top.scala 490:26:@660.28]
  assign _T_596 = $signed(wx) + $signed(_T_594); // @[collide_top.scala 490:26:@661.28]
  assign _T_597 = $signed(_T_596); // @[collide_top.scala 490:26:@662.28]
  assign _T_598 = tcvx[14:6]; // @[collide_top.scala 490:52:@663.28]
  assign _T_599 = $signed(_T_598); // @[collide_top.scala 490:59:@664.28]
  assign _T_600 = $signed(_T_597) - $signed(_T_599); // @[collide_top.scala 490:46:@665.28]
  assign _T_601 = $signed(_T_597) - $signed(_T_599); // @[collide_top.scala 490:46:@666.28]
  assign _T_602 = $signed(_T_601); // @[collide_top.scala 490:46:@667.28]
  assign _T_603 = scuy[14:6]; // @[collide_top.scala 491:32:@669.28]
  assign _T_604 = $signed(_T_603); // @[collide_top.scala 491:39:@670.28]
  assign _T_605 = $signed(wy) + $signed(_T_604); // @[collide_top.scala 491:26:@671.28]
  assign _T_606 = $signed(wy) + $signed(_T_604); // @[collide_top.scala 491:26:@672.28]
  assign _T_607 = $signed(_T_606); // @[collide_top.scala 491:26:@673.28]
  assign _T_608 = tcvy[14:6]; // @[collide_top.scala 491:52:@674.28]
  assign _T_609 = $signed(_T_608); // @[collide_top.scala 491:59:@675.28]
  assign _T_610 = $signed(_T_607) - $signed(_T_609); // @[collide_top.scala 491:46:@676.28]
  assign _T_611 = $signed(_T_607) - $signed(_T_609); // @[collide_top.scala 491:46:@677.28]
  assign _T_612 = $signed(_T_611); // @[collide_top.scala 491:46:@678.28]
  assign _T_613 = scuz[14:6]; // @[collide_top.scala 492:32:@680.28]
  assign _T_614 = $signed(_T_613); // @[collide_top.scala 492:39:@681.28]
  assign _T_615 = $signed(wz) + $signed(_T_614); // @[collide_top.scala 492:26:@682.28]
  assign _T_616 = $signed(wz) + $signed(_T_614); // @[collide_top.scala 492:26:@683.28]
  assign _T_617 = $signed(_T_616); // @[collide_top.scala 492:26:@684.28]
  assign _T_618 = tcvz[14:6]; // @[collide_top.scala 492:52:@685.28]
  assign _T_619 = $signed(_T_618); // @[collide_top.scala 492:59:@686.28]
  assign _T_620 = $signed(_T_617) - $signed(_T_619); // @[collide_top.scala 492:46:@687.28]
  assign _T_621 = $signed(_T_617) - $signed(_T_619); // @[collide_top.scala 492:46:@688.28]
  assign _T_622 = $signed(_T_621); // @[collide_top.scala 492:46:@689.28]
  assign _T_624 = io_state == 8'h16; // @[collide_top.scala 494:29:@693.28]
  assign _T_625 = $signed(dx) * $signed(dx); // @[collide_top.scala 496:28:@695.30]
  assign _T_626 = $signed(dy) * $signed(dy); // @[collide_top.scala 497:28:@697.30]
  assign _T_627 = $signed(dz) * $signed(dz); // @[collide_top.scala 498:28:@699.30]
  assign _T_629 = io_state == 8'h17; // @[collide_top.scala 500:29:@703.30]
  assign _T_630 = $signed(dxdx) + $signed(dydy); // @[collide_top.scala 502:38:@705.32]
  assign _T_631 = $signed(dxdx) + $signed(dydy); // @[collide_top.scala 502:38:@706.32]
  assign _T_632 = $signed(_T_631); // @[collide_top.scala 502:38:@707.32]
  assign _T_633 = $signed(_T_632) + $signed(dzdz); // @[collide_top.scala 502:45:@708.32]
  assign _T_634 = $signed(_T_632) + $signed(dzdz); // @[collide_top.scala 502:45:@709.32]
  assign _T_635 = $signed(_T_634); // @[collide_top.scala 502:45:@710.32]
  assign _T_637 = io_state == 8'h18; // @[collide_top.scala 504:29:@714.32]
  assign _GEN_0 = _T_637 ? $signed(_T_635) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_1 = _T_637 ? $signed(ux) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_2 = _T_637 ? $signed(uy) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_3 = _T_637 ? $signed(uz) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_4 = _T_637 ? $signed(vx) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_5 = _T_637 ? $signed(vy) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_6 = _T_637 ? $signed(vz) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_7 = _T_637 ? $signed(wx) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_8 = _T_637 ? $signed(wy) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_9 = _T_637 ? $signed(wz) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_10 = _T_637 ? $signed(uxux) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_11 = _T_637 ? $signed(uyuy) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_12 = _T_637 ? $signed(uzuz) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_13 = _T_637 ? $signed(uxvx) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_14 = _T_637 ? $signed(uyvy) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_15 = _T_637 ? $signed(uzvz) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_16 = _T_637 ? $signed(vxvx) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_17 = _T_637 ? $signed(vyvy) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_18 = _T_637 ? $signed(vzvz) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_19 = _T_637 ? $signed(uxwx) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_20 = _T_637 ? $signed(uywy) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_21 = _T_637 ? $signed(uzwz) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_22 = _T_637 ? $signed(vxwx) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_23 = _T_637 ? $signed(vywy) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_24 = _T_637 ? $signed(vzwz) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_25 = _T_637 ? $signed(a) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_26 = _T_637 ? $signed(b) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_27 = _T_637 ? $signed(c) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_28 = _T_637 ? $signed(d) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_29 = _T_637 ? $signed(e) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_30 = _T_637 ? $signed(a_ex) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_31 = _T_637 ? $signed(b_ex) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_32 = _T_637 ? $signed(c_ex) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_33 = _T_637 ? $signed(d_ex) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_34 = _T_637 ? $signed(e_ex) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_35 = _T_637 ? $signed(ac) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_36 = _T_637 ? $signed(bb) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_37 = _T_637 ? $signed(be) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_38 = _T_637 ? $signed(cd) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_39 = _T_637 ? $signed(ae) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_40 = _T_637 ? $signed(bd) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_41 = _T_637 ? $signed(D_SUB_B) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_42 = _T_637 ? $signed(sn_temp) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_43 = _T_637 ? $signed(sd_temp) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_44 = _T_637 ? $signed(tn_temp) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_45 = _T_637 ? $signed(td) : $signed(36'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_46 = _T_637 ? sc : 6'h0; // @[collide_top.scala 505:9:@715.32]
  assign _GEN_47 = _T_637 ? tc : 6'h0; // @[collide_top.scala 505:9:@715.32]
  assign _GEN_48 = _T_637 ? sn_calData : 41'h0; // @[collide_top.scala 505:9:@715.32]
  assign _GEN_49 = _T_637 ? sd_calData : 41'h0; // @[collide_top.scala 505:9:@715.32]
  assign _GEN_50 = _T_637 ? td_calData : 41'h0; // @[collide_top.scala 505:9:@715.32]
  assign _GEN_51 = _T_637 ? $signed(scux) : $signed(15'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_52 = _T_637 ? $signed(tcvx) : $signed(15'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_53 = _T_637 ? $signed(scuy) : $signed(15'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_54 = _T_637 ? $signed(tcvy) : $signed(15'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_55 = _T_637 ? $signed(scuz) : $signed(15'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_56 = _T_637 ? $signed(tcvz) : $signed(15'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_57 = _T_637 ? $signed(dx) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_58 = _T_637 ? $signed(dy) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_59 = _T_637 ? $signed(dz) : $signed(9'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_60 = _T_637 ? $signed(dxdx) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_61 = _T_637 ? $signed(dydy) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_62 = _T_637 ? $signed(dzdz) : $signed(18'sh0); // @[collide_top.scala 505:9:@715.32]
  assign _GEN_63 = _T_629 ? $signed(_T_635) : $signed(_GEN_0); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_64 = _T_629 ? $signed(ux) : $signed(_GEN_1); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_65 = _T_629 ? $signed(uy) : $signed(_GEN_2); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_66 = _T_629 ? $signed(uz) : $signed(_GEN_3); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_67 = _T_629 ? $signed(vx) : $signed(_GEN_4); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_68 = _T_629 ? $signed(vy) : $signed(_GEN_5); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_69 = _T_629 ? $signed(vz) : $signed(_GEN_6); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_70 = _T_629 ? $signed(wx) : $signed(_GEN_7); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_71 = _T_629 ? $signed(wy) : $signed(_GEN_8); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_72 = _T_629 ? $signed(wz) : $signed(_GEN_9); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_73 = _T_629 ? $signed(uxux) : $signed(_GEN_10); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_74 = _T_629 ? $signed(uyuy) : $signed(_GEN_11); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_75 = _T_629 ? $signed(uzuz) : $signed(_GEN_12); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_76 = _T_629 ? $signed(uxvx) : $signed(_GEN_13); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_77 = _T_629 ? $signed(uyvy) : $signed(_GEN_14); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_78 = _T_629 ? $signed(uzvz) : $signed(_GEN_15); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_79 = _T_629 ? $signed(vxvx) : $signed(_GEN_16); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_80 = _T_629 ? $signed(vyvy) : $signed(_GEN_17); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_81 = _T_629 ? $signed(vzvz) : $signed(_GEN_18); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_82 = _T_629 ? $signed(uxwx) : $signed(_GEN_19); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_83 = _T_629 ? $signed(uywy) : $signed(_GEN_20); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_84 = _T_629 ? $signed(uzwz) : $signed(_GEN_21); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_85 = _T_629 ? $signed(vxwx) : $signed(_GEN_22); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_86 = _T_629 ? $signed(vywy) : $signed(_GEN_23); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_87 = _T_629 ? $signed(vzwz) : $signed(_GEN_24); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_88 = _T_629 ? $signed(a) : $signed(_GEN_25); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_89 = _T_629 ? $signed(b) : $signed(_GEN_26); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_90 = _T_629 ? $signed(c) : $signed(_GEN_27); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_91 = _T_629 ? $signed(d) : $signed(_GEN_28); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_92 = _T_629 ? $signed(e) : $signed(_GEN_29); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_93 = _T_629 ? $signed(a_ex) : $signed(_GEN_30); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_94 = _T_629 ? $signed(b_ex) : $signed(_GEN_31); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_95 = _T_629 ? $signed(c_ex) : $signed(_GEN_32); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_96 = _T_629 ? $signed(d_ex) : $signed(_GEN_33); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_97 = _T_629 ? $signed(e_ex) : $signed(_GEN_34); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_98 = _T_629 ? $signed(ac) : $signed(_GEN_35); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_99 = _T_629 ? $signed(bb) : $signed(_GEN_36); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_100 = _T_629 ? $signed(be) : $signed(_GEN_37); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_101 = _T_629 ? $signed(cd) : $signed(_GEN_38); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_102 = _T_629 ? $signed(ae) : $signed(_GEN_39); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_103 = _T_629 ? $signed(bd) : $signed(_GEN_40); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_104 = _T_629 ? $signed(D_SUB_B) : $signed(_GEN_41); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_105 = _T_629 ? $signed(sn_temp) : $signed(_GEN_42); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_106 = _T_629 ? $signed(sd_temp) : $signed(_GEN_43); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_107 = _T_629 ? $signed(tn_temp) : $signed(_GEN_44); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_108 = _T_629 ? $signed(td) : $signed(_GEN_45); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_109 = _T_629 ? sc : _GEN_46; // @[collide_top.scala 501:9:@704.30]
  assign _GEN_110 = _T_629 ? tc : _GEN_47; // @[collide_top.scala 501:9:@704.30]
  assign _GEN_111 = _T_629 ? sn_calData : _GEN_48; // @[collide_top.scala 501:9:@704.30]
  assign _GEN_112 = _T_629 ? sd_calData : _GEN_49; // @[collide_top.scala 501:9:@704.30]
  assign _GEN_113 = _T_629 ? td_calData : _GEN_50; // @[collide_top.scala 501:9:@704.30]
  assign _GEN_114 = _T_629 ? $signed(scux) : $signed(_GEN_51); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_115 = _T_629 ? $signed(tcvx) : $signed(_GEN_52); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_116 = _T_629 ? $signed(scuy) : $signed(_GEN_53); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_117 = _T_629 ? $signed(tcvy) : $signed(_GEN_54); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_118 = _T_629 ? $signed(scuz) : $signed(_GEN_55); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_119 = _T_629 ? $signed(tcvz) : $signed(_GEN_56); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_120 = _T_629 ? $signed(dx) : $signed(_GEN_57); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_121 = _T_629 ? $signed(dy) : $signed(_GEN_58); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_122 = _T_629 ? $signed(dz) : $signed(_GEN_59); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_123 = _T_629 ? $signed(dxdx) : $signed(_GEN_60); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_124 = _T_629 ? $signed(dydy) : $signed(_GEN_61); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_125 = _T_629 ? $signed(dzdz) : $signed(_GEN_62); // @[collide_top.scala 501:9:@704.30]
  assign _GEN_126 = _T_624 ? $signed(_T_625) : $signed(_GEN_123); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_127 = _T_624 ? $signed(_T_626) : $signed(_GEN_124); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_128 = _T_624 ? $signed(_T_627) : $signed(_GEN_125); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_129 = _T_624 ? $signed(distance_Reg) : $signed(_GEN_63); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_130 = _T_624 ? $signed(ux) : $signed(_GEN_64); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_131 = _T_624 ? $signed(uy) : $signed(_GEN_65); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_132 = _T_624 ? $signed(uz) : $signed(_GEN_66); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_133 = _T_624 ? $signed(vx) : $signed(_GEN_67); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_134 = _T_624 ? $signed(vy) : $signed(_GEN_68); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_135 = _T_624 ? $signed(vz) : $signed(_GEN_69); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_136 = _T_624 ? $signed(wx) : $signed(_GEN_70); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_137 = _T_624 ? $signed(wy) : $signed(_GEN_71); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_138 = _T_624 ? $signed(wz) : $signed(_GEN_72); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_139 = _T_624 ? $signed(uxux) : $signed(_GEN_73); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_140 = _T_624 ? $signed(uyuy) : $signed(_GEN_74); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_141 = _T_624 ? $signed(uzuz) : $signed(_GEN_75); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_142 = _T_624 ? $signed(uxvx) : $signed(_GEN_76); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_143 = _T_624 ? $signed(uyvy) : $signed(_GEN_77); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_144 = _T_624 ? $signed(uzvz) : $signed(_GEN_78); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_145 = _T_624 ? $signed(vxvx) : $signed(_GEN_79); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_146 = _T_624 ? $signed(vyvy) : $signed(_GEN_80); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_147 = _T_624 ? $signed(vzvz) : $signed(_GEN_81); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_148 = _T_624 ? $signed(uxwx) : $signed(_GEN_82); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_149 = _T_624 ? $signed(uywy) : $signed(_GEN_83); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_150 = _T_624 ? $signed(uzwz) : $signed(_GEN_84); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_151 = _T_624 ? $signed(vxwx) : $signed(_GEN_85); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_152 = _T_624 ? $signed(vywy) : $signed(_GEN_86); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_153 = _T_624 ? $signed(vzwz) : $signed(_GEN_87); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_154 = _T_624 ? $signed(a) : $signed(_GEN_88); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_155 = _T_624 ? $signed(b) : $signed(_GEN_89); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_156 = _T_624 ? $signed(c) : $signed(_GEN_90); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_157 = _T_624 ? $signed(d) : $signed(_GEN_91); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_158 = _T_624 ? $signed(e) : $signed(_GEN_92); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_159 = _T_624 ? $signed(a_ex) : $signed(_GEN_93); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_160 = _T_624 ? $signed(b_ex) : $signed(_GEN_94); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_161 = _T_624 ? $signed(c_ex) : $signed(_GEN_95); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_162 = _T_624 ? $signed(d_ex) : $signed(_GEN_96); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_163 = _T_624 ? $signed(e_ex) : $signed(_GEN_97); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_164 = _T_624 ? $signed(ac) : $signed(_GEN_98); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_165 = _T_624 ? $signed(bb) : $signed(_GEN_99); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_166 = _T_624 ? $signed(be) : $signed(_GEN_100); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_167 = _T_624 ? $signed(cd) : $signed(_GEN_101); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_168 = _T_624 ? $signed(ae) : $signed(_GEN_102); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_169 = _T_624 ? $signed(bd) : $signed(_GEN_103); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_170 = _T_624 ? $signed(D_SUB_B) : $signed(_GEN_104); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_171 = _T_624 ? $signed(sn_temp) : $signed(_GEN_105); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_172 = _T_624 ? $signed(sd_temp) : $signed(_GEN_106); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_173 = _T_624 ? $signed(tn_temp) : $signed(_GEN_107); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_174 = _T_624 ? $signed(td) : $signed(_GEN_108); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_175 = _T_624 ? sc : _GEN_109; // @[collide_top.scala 495:9:@694.28]
  assign _GEN_176 = _T_624 ? tc : _GEN_110; // @[collide_top.scala 495:9:@694.28]
  assign _GEN_177 = _T_624 ? sn_calData : _GEN_111; // @[collide_top.scala 495:9:@694.28]
  assign _GEN_178 = _T_624 ? sd_calData : _GEN_112; // @[collide_top.scala 495:9:@694.28]
  assign _GEN_179 = _T_624 ? td_calData : _GEN_113; // @[collide_top.scala 495:9:@694.28]
  assign _GEN_180 = _T_624 ? $signed(scux) : $signed(_GEN_114); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_181 = _T_624 ? $signed(tcvx) : $signed(_GEN_115); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_182 = _T_624 ? $signed(scuy) : $signed(_GEN_116); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_183 = _T_624 ? $signed(tcvy) : $signed(_GEN_117); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_184 = _T_624 ? $signed(scuz) : $signed(_GEN_118); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_185 = _T_624 ? $signed(tcvz) : $signed(_GEN_119); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_186 = _T_624 ? $signed(dx) : $signed(_GEN_120); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_187 = _T_624 ? $signed(dy) : $signed(_GEN_121); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_188 = _T_624 ? $signed(dz) : $signed(_GEN_122); // @[collide_top.scala 495:9:@694.28]
  assign _GEN_189 = _T_592 ? $signed(_T_602) : $signed(_GEN_186); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_190 = _T_592 ? $signed(_T_612) : $signed(_GEN_187); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_191 = _T_592 ? $signed(_T_622) : $signed(_GEN_188); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_192 = _T_592 ? $signed(dxdx) : $signed(_GEN_126); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_193 = _T_592 ? $signed(dydy) : $signed(_GEN_127); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_194 = _T_592 ? $signed(dzdz) : $signed(_GEN_128); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_195 = _T_592 ? $signed(distance_Reg) : $signed(_GEN_129); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_196 = _T_592 ? $signed(ux) : $signed(_GEN_130); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_197 = _T_592 ? $signed(uy) : $signed(_GEN_131); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_198 = _T_592 ? $signed(uz) : $signed(_GEN_132); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_199 = _T_592 ? $signed(vx) : $signed(_GEN_133); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_200 = _T_592 ? $signed(vy) : $signed(_GEN_134); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_201 = _T_592 ? $signed(vz) : $signed(_GEN_135); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_202 = _T_592 ? $signed(wx) : $signed(_GEN_136); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_203 = _T_592 ? $signed(wy) : $signed(_GEN_137); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_204 = _T_592 ? $signed(wz) : $signed(_GEN_138); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_205 = _T_592 ? $signed(uxux) : $signed(_GEN_139); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_206 = _T_592 ? $signed(uyuy) : $signed(_GEN_140); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_207 = _T_592 ? $signed(uzuz) : $signed(_GEN_141); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_208 = _T_592 ? $signed(uxvx) : $signed(_GEN_142); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_209 = _T_592 ? $signed(uyvy) : $signed(_GEN_143); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_210 = _T_592 ? $signed(uzvz) : $signed(_GEN_144); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_211 = _T_592 ? $signed(vxvx) : $signed(_GEN_145); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_212 = _T_592 ? $signed(vyvy) : $signed(_GEN_146); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_213 = _T_592 ? $signed(vzvz) : $signed(_GEN_147); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_214 = _T_592 ? $signed(uxwx) : $signed(_GEN_148); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_215 = _T_592 ? $signed(uywy) : $signed(_GEN_149); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_216 = _T_592 ? $signed(uzwz) : $signed(_GEN_150); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_217 = _T_592 ? $signed(vxwx) : $signed(_GEN_151); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_218 = _T_592 ? $signed(vywy) : $signed(_GEN_152); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_219 = _T_592 ? $signed(vzwz) : $signed(_GEN_153); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_220 = _T_592 ? $signed(a) : $signed(_GEN_154); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_221 = _T_592 ? $signed(b) : $signed(_GEN_155); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_222 = _T_592 ? $signed(c) : $signed(_GEN_156); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_223 = _T_592 ? $signed(d) : $signed(_GEN_157); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_224 = _T_592 ? $signed(e) : $signed(_GEN_158); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_225 = _T_592 ? $signed(a_ex) : $signed(_GEN_159); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_226 = _T_592 ? $signed(b_ex) : $signed(_GEN_160); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_227 = _T_592 ? $signed(c_ex) : $signed(_GEN_161); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_228 = _T_592 ? $signed(d_ex) : $signed(_GEN_162); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_229 = _T_592 ? $signed(e_ex) : $signed(_GEN_163); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_230 = _T_592 ? $signed(ac) : $signed(_GEN_164); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_231 = _T_592 ? $signed(bb) : $signed(_GEN_165); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_232 = _T_592 ? $signed(be) : $signed(_GEN_166); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_233 = _T_592 ? $signed(cd) : $signed(_GEN_167); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_234 = _T_592 ? $signed(ae) : $signed(_GEN_168); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_235 = _T_592 ? $signed(bd) : $signed(_GEN_169); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_236 = _T_592 ? $signed(D_SUB_B) : $signed(_GEN_170); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_237 = _T_592 ? $signed(sn_temp) : $signed(_GEN_171); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_238 = _T_592 ? $signed(sd_temp) : $signed(_GEN_172); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_239 = _T_592 ? $signed(tn_temp) : $signed(_GEN_173); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_240 = _T_592 ? $signed(td) : $signed(_GEN_174); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_241 = _T_592 ? sc : _GEN_175; // @[collide_top.scala 489:9:@657.26]
  assign _GEN_242 = _T_592 ? tc : _GEN_176; // @[collide_top.scala 489:9:@657.26]
  assign _GEN_243 = _T_592 ? sn_calData : _GEN_177; // @[collide_top.scala 489:9:@657.26]
  assign _GEN_244 = _T_592 ? sd_calData : _GEN_178; // @[collide_top.scala 489:9:@657.26]
  assign _GEN_245 = _T_592 ? td_calData : _GEN_179; // @[collide_top.scala 489:9:@657.26]
  assign _GEN_246 = _T_592 ? $signed(scux) : $signed(_GEN_180); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_247 = _T_592 ? $signed(tcvx) : $signed(_GEN_181); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_248 = _T_592 ? $signed(scuy) : $signed(_GEN_182); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_249 = _T_592 ? $signed(tcvy) : $signed(_GEN_183); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_250 = _T_592 ? $signed(scuz) : $signed(_GEN_184); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_251 = _T_592 ? $signed(tcvz) : $signed(_GEN_185); // @[collide_top.scala 489:9:@657.26]
  assign _GEN_252 = _T_566 ? $signed(_T_570) : $signed(_GEN_246); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_253 = _T_566 ? $signed(_T_574) : $signed(_GEN_247); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_254 = _T_566 ? $signed(_T_578) : $signed(_GEN_248); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_255 = _T_566 ? $signed(_T_582) : $signed(_GEN_249); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_256 = _T_566 ? $signed(_T_586) : $signed(_GEN_250); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_257 = _T_566 ? $signed(_T_590) : $signed(_GEN_251); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_258 = _T_566 ? $signed(dx) : $signed(_GEN_189); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_259 = _T_566 ? $signed(dy) : $signed(_GEN_190); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_260 = _T_566 ? $signed(dz) : $signed(_GEN_191); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_261 = _T_566 ? $signed(dxdx) : $signed(_GEN_192); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_262 = _T_566 ? $signed(dydy) : $signed(_GEN_193); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_263 = _T_566 ? $signed(dzdz) : $signed(_GEN_194); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_264 = _T_566 ? $signed(distance_Reg) : $signed(_GEN_195); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_265 = _T_566 ? $signed(ux) : $signed(_GEN_196); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_266 = _T_566 ? $signed(uy) : $signed(_GEN_197); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_267 = _T_566 ? $signed(uz) : $signed(_GEN_198); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_268 = _T_566 ? $signed(vx) : $signed(_GEN_199); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_269 = _T_566 ? $signed(vy) : $signed(_GEN_200); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_270 = _T_566 ? $signed(vz) : $signed(_GEN_201); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_271 = _T_566 ? $signed(wx) : $signed(_GEN_202); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_272 = _T_566 ? $signed(wy) : $signed(_GEN_203); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_273 = _T_566 ? $signed(wz) : $signed(_GEN_204); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_274 = _T_566 ? $signed(uxux) : $signed(_GEN_205); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_275 = _T_566 ? $signed(uyuy) : $signed(_GEN_206); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_276 = _T_566 ? $signed(uzuz) : $signed(_GEN_207); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_277 = _T_566 ? $signed(uxvx) : $signed(_GEN_208); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_278 = _T_566 ? $signed(uyvy) : $signed(_GEN_209); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_279 = _T_566 ? $signed(uzvz) : $signed(_GEN_210); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_280 = _T_566 ? $signed(vxvx) : $signed(_GEN_211); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_281 = _T_566 ? $signed(vyvy) : $signed(_GEN_212); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_282 = _T_566 ? $signed(vzvz) : $signed(_GEN_213); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_283 = _T_566 ? $signed(uxwx) : $signed(_GEN_214); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_284 = _T_566 ? $signed(uywy) : $signed(_GEN_215); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_285 = _T_566 ? $signed(uzwz) : $signed(_GEN_216); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_286 = _T_566 ? $signed(vxwx) : $signed(_GEN_217); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_287 = _T_566 ? $signed(vywy) : $signed(_GEN_218); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_288 = _T_566 ? $signed(vzwz) : $signed(_GEN_219); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_289 = _T_566 ? $signed(a) : $signed(_GEN_220); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_290 = _T_566 ? $signed(b) : $signed(_GEN_221); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_291 = _T_566 ? $signed(c) : $signed(_GEN_222); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_292 = _T_566 ? $signed(d) : $signed(_GEN_223); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_293 = _T_566 ? $signed(e) : $signed(_GEN_224); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_294 = _T_566 ? $signed(a_ex) : $signed(_GEN_225); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_295 = _T_566 ? $signed(b_ex) : $signed(_GEN_226); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_296 = _T_566 ? $signed(c_ex) : $signed(_GEN_227); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_297 = _T_566 ? $signed(d_ex) : $signed(_GEN_228); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_298 = _T_566 ? $signed(e_ex) : $signed(_GEN_229); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_299 = _T_566 ? $signed(ac) : $signed(_GEN_230); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_300 = _T_566 ? $signed(bb) : $signed(_GEN_231); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_301 = _T_566 ? $signed(be) : $signed(_GEN_232); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_302 = _T_566 ? $signed(cd) : $signed(_GEN_233); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_303 = _T_566 ? $signed(ae) : $signed(_GEN_234); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_304 = _T_566 ? $signed(bd) : $signed(_GEN_235); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_305 = _T_566 ? $signed(D_SUB_B) : $signed(_GEN_236); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_306 = _T_566 ? $signed(sn_temp) : $signed(_GEN_237); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_307 = _T_566 ? $signed(sd_temp) : $signed(_GEN_238); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_308 = _T_566 ? $signed(tn_temp) : $signed(_GEN_239); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_309 = _T_566 ? $signed(td) : $signed(_GEN_240); // @[collide_top.scala 480:9:@623.24]
  assign _GEN_310 = _T_566 ? sc : _GEN_241; // @[collide_top.scala 480:9:@623.24]
  assign _GEN_311 = _T_566 ? tc : _GEN_242; // @[collide_top.scala 480:9:@623.24]
  assign _GEN_312 = _T_566 ? sn_calData : _GEN_243; // @[collide_top.scala 480:9:@623.24]
  assign _GEN_313 = _T_566 ? sd_calData : _GEN_244; // @[collide_top.scala 480:9:@623.24]
  assign _GEN_314 = _T_566 ? td_calData : _GEN_245; // @[collide_top.scala 480:9:@623.24]
  assign _GEN_315 = _T_544 ? _T_504 : _GEN_312; // @[collide_top.scala 472:9:@597.22]
  assign _GEN_316 = _T_544 ? _T_510 : {{1'd0}, _GEN_310}; // @[collide_top.scala 472:9:@597.22]
  assign _GEN_317 = _T_544 ? _T_514 : tn_calData; // @[collide_top.scala 472:9:@597.22]
  assign _GEN_318 = _T_544 ? _T_520 : {{1'd0}, _GEN_311}; // @[collide_top.scala 472:9:@597.22]
  assign _GEN_319 = _T_544 ? $signed(scux) : $signed(_GEN_252); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_320 = _T_544 ? $signed(tcvx) : $signed(_GEN_253); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_321 = _T_544 ? $signed(scuy) : $signed(_GEN_254); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_322 = _T_544 ? $signed(tcvy) : $signed(_GEN_255); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_323 = _T_544 ? $signed(scuz) : $signed(_GEN_256); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_324 = _T_544 ? $signed(tcvz) : $signed(_GEN_257); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_325 = _T_544 ? $signed(dx) : $signed(_GEN_258); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_326 = _T_544 ? $signed(dy) : $signed(_GEN_259); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_327 = _T_544 ? $signed(dz) : $signed(_GEN_260); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_328 = _T_544 ? $signed(dxdx) : $signed(_GEN_261); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_329 = _T_544 ? $signed(dydy) : $signed(_GEN_262); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_330 = _T_544 ? $signed(dzdz) : $signed(_GEN_263); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_331 = _T_544 ? $signed(distance_Reg) : $signed(_GEN_264); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_332 = _T_544 ? $signed(ux) : $signed(_GEN_265); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_333 = _T_544 ? $signed(uy) : $signed(_GEN_266); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_334 = _T_544 ? $signed(uz) : $signed(_GEN_267); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_335 = _T_544 ? $signed(vx) : $signed(_GEN_268); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_336 = _T_544 ? $signed(vy) : $signed(_GEN_269); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_337 = _T_544 ? $signed(vz) : $signed(_GEN_270); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_338 = _T_544 ? $signed(wx) : $signed(_GEN_271); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_339 = _T_544 ? $signed(wy) : $signed(_GEN_272); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_340 = _T_544 ? $signed(wz) : $signed(_GEN_273); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_341 = _T_544 ? $signed(uxux) : $signed(_GEN_274); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_342 = _T_544 ? $signed(uyuy) : $signed(_GEN_275); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_343 = _T_544 ? $signed(uzuz) : $signed(_GEN_276); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_344 = _T_544 ? $signed(uxvx) : $signed(_GEN_277); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_345 = _T_544 ? $signed(uyvy) : $signed(_GEN_278); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_346 = _T_544 ? $signed(uzvz) : $signed(_GEN_279); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_347 = _T_544 ? $signed(vxvx) : $signed(_GEN_280); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_348 = _T_544 ? $signed(vyvy) : $signed(_GEN_281); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_349 = _T_544 ? $signed(vzvz) : $signed(_GEN_282); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_350 = _T_544 ? $signed(uxwx) : $signed(_GEN_283); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_351 = _T_544 ? $signed(uywy) : $signed(_GEN_284); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_352 = _T_544 ? $signed(uzwz) : $signed(_GEN_285); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_353 = _T_544 ? $signed(vxwx) : $signed(_GEN_286); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_354 = _T_544 ? $signed(vywy) : $signed(_GEN_287); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_355 = _T_544 ? $signed(vzwz) : $signed(_GEN_288); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_356 = _T_544 ? $signed(a) : $signed(_GEN_289); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_357 = _T_544 ? $signed(b) : $signed(_GEN_290); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_358 = _T_544 ? $signed(c) : $signed(_GEN_291); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_359 = _T_544 ? $signed(d) : $signed(_GEN_292); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_360 = _T_544 ? $signed(e) : $signed(_GEN_293); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_361 = _T_544 ? $signed(a_ex) : $signed(_GEN_294); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_362 = _T_544 ? $signed(b_ex) : $signed(_GEN_295); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_363 = _T_544 ? $signed(c_ex) : $signed(_GEN_296); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_364 = _T_544 ? $signed(d_ex) : $signed(_GEN_297); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_365 = _T_544 ? $signed(e_ex) : $signed(_GEN_298); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_366 = _T_544 ? $signed(ac) : $signed(_GEN_299); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_367 = _T_544 ? $signed(bb) : $signed(_GEN_300); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_368 = _T_544 ? $signed(be) : $signed(_GEN_301); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_369 = _T_544 ? $signed(cd) : $signed(_GEN_302); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_370 = _T_544 ? $signed(ae) : $signed(_GEN_303); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_371 = _T_544 ? $signed(bd) : $signed(_GEN_304); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_372 = _T_544 ? $signed(D_SUB_B) : $signed(_GEN_305); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_373 = _T_544 ? $signed(sn_temp) : $signed(_GEN_306); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_374 = _T_544 ? $signed(sd_temp) : $signed(_GEN_307); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_375 = _T_544 ? $signed(tn_temp) : $signed(_GEN_308); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_376 = _T_544 ? $signed(td) : $signed(_GEN_309); // @[collide_top.scala 472:9:@597.22]
  assign _GEN_377 = _T_544 ? sd_calData : _GEN_313; // @[collide_top.scala 472:9:@597.22]
  assign _GEN_378 = _T_544 ? td_calData : _GEN_314; // @[collide_top.scala 472:9:@597.22]
  assign _GEN_379 = _T_522 ? _T_504 : _GEN_315; // @[collide_top.scala 464:9:@571.20]
  assign _GEN_380 = _T_522 ? _T_510 : _GEN_316; // @[collide_top.scala 464:9:@571.20]
  assign _GEN_381 = _T_522 ? _T_514 : _GEN_317; // @[collide_top.scala 464:9:@571.20]
  assign _GEN_382 = _T_522 ? _T_520 : _GEN_318; // @[collide_top.scala 464:9:@571.20]
  assign _GEN_383 = _T_522 ? $signed(scux) : $signed(_GEN_319); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_384 = _T_522 ? $signed(tcvx) : $signed(_GEN_320); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_385 = _T_522 ? $signed(scuy) : $signed(_GEN_321); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_386 = _T_522 ? $signed(tcvy) : $signed(_GEN_322); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_387 = _T_522 ? $signed(scuz) : $signed(_GEN_323); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_388 = _T_522 ? $signed(tcvz) : $signed(_GEN_324); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_389 = _T_522 ? $signed(dx) : $signed(_GEN_325); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_390 = _T_522 ? $signed(dy) : $signed(_GEN_326); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_391 = _T_522 ? $signed(dz) : $signed(_GEN_327); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_392 = _T_522 ? $signed(dxdx) : $signed(_GEN_328); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_393 = _T_522 ? $signed(dydy) : $signed(_GEN_329); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_394 = _T_522 ? $signed(dzdz) : $signed(_GEN_330); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_395 = _T_522 ? $signed(distance_Reg) : $signed(_GEN_331); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_396 = _T_522 ? $signed(ux) : $signed(_GEN_332); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_397 = _T_522 ? $signed(uy) : $signed(_GEN_333); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_398 = _T_522 ? $signed(uz) : $signed(_GEN_334); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_399 = _T_522 ? $signed(vx) : $signed(_GEN_335); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_400 = _T_522 ? $signed(vy) : $signed(_GEN_336); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_401 = _T_522 ? $signed(vz) : $signed(_GEN_337); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_402 = _T_522 ? $signed(wx) : $signed(_GEN_338); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_403 = _T_522 ? $signed(wy) : $signed(_GEN_339); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_404 = _T_522 ? $signed(wz) : $signed(_GEN_340); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_405 = _T_522 ? $signed(uxux) : $signed(_GEN_341); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_406 = _T_522 ? $signed(uyuy) : $signed(_GEN_342); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_407 = _T_522 ? $signed(uzuz) : $signed(_GEN_343); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_408 = _T_522 ? $signed(uxvx) : $signed(_GEN_344); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_409 = _T_522 ? $signed(uyvy) : $signed(_GEN_345); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_410 = _T_522 ? $signed(uzvz) : $signed(_GEN_346); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_411 = _T_522 ? $signed(vxvx) : $signed(_GEN_347); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_412 = _T_522 ? $signed(vyvy) : $signed(_GEN_348); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_413 = _T_522 ? $signed(vzvz) : $signed(_GEN_349); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_414 = _T_522 ? $signed(uxwx) : $signed(_GEN_350); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_415 = _T_522 ? $signed(uywy) : $signed(_GEN_351); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_416 = _T_522 ? $signed(uzwz) : $signed(_GEN_352); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_417 = _T_522 ? $signed(vxwx) : $signed(_GEN_353); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_418 = _T_522 ? $signed(vywy) : $signed(_GEN_354); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_419 = _T_522 ? $signed(vzwz) : $signed(_GEN_355); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_420 = _T_522 ? $signed(a) : $signed(_GEN_356); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_421 = _T_522 ? $signed(b) : $signed(_GEN_357); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_422 = _T_522 ? $signed(c) : $signed(_GEN_358); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_423 = _T_522 ? $signed(d) : $signed(_GEN_359); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_424 = _T_522 ? $signed(e) : $signed(_GEN_360); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_425 = _T_522 ? $signed(a_ex) : $signed(_GEN_361); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_426 = _T_522 ? $signed(b_ex) : $signed(_GEN_362); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_427 = _T_522 ? $signed(c_ex) : $signed(_GEN_363); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_428 = _T_522 ? $signed(d_ex) : $signed(_GEN_364); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_429 = _T_522 ? $signed(e_ex) : $signed(_GEN_365); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_430 = _T_522 ? $signed(ac) : $signed(_GEN_366); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_431 = _T_522 ? $signed(bb) : $signed(_GEN_367); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_432 = _T_522 ? $signed(be) : $signed(_GEN_368); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_433 = _T_522 ? $signed(cd) : $signed(_GEN_369); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_434 = _T_522 ? $signed(ae) : $signed(_GEN_370); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_435 = _T_522 ? $signed(bd) : $signed(_GEN_371); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_436 = _T_522 ? $signed(D_SUB_B) : $signed(_GEN_372); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_437 = _T_522 ? $signed(sn_temp) : $signed(_GEN_373); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_438 = _T_522 ? $signed(sd_temp) : $signed(_GEN_374); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_439 = _T_522 ? $signed(tn_temp) : $signed(_GEN_375); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_440 = _T_522 ? $signed(td) : $signed(_GEN_376); // @[collide_top.scala 464:9:@571.20]
  assign _GEN_441 = _T_522 ? sd_calData : _GEN_377; // @[collide_top.scala 464:9:@571.20]
  assign _GEN_442 = _T_522 ? td_calData : _GEN_378; // @[collide_top.scala 464:9:@571.20]
  assign _GEN_443 = _T_500 ? _T_504 : _GEN_379; // @[collide_top.scala 455:9:@545.18]
  assign _GEN_444 = _T_500 ? _T_510 : _GEN_380; // @[collide_top.scala 455:9:@545.18]
  assign _GEN_445 = _T_500 ? _T_514 : _GEN_381; // @[collide_top.scala 455:9:@545.18]
  assign _GEN_446 = _T_500 ? _T_520 : _GEN_382; // @[collide_top.scala 455:9:@545.18]
  assign _GEN_447 = _T_500 ? $signed(scux) : $signed(_GEN_383); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_448 = _T_500 ? $signed(tcvx) : $signed(_GEN_384); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_449 = _T_500 ? $signed(scuy) : $signed(_GEN_385); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_450 = _T_500 ? $signed(tcvy) : $signed(_GEN_386); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_451 = _T_500 ? $signed(scuz) : $signed(_GEN_387); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_452 = _T_500 ? $signed(tcvz) : $signed(_GEN_388); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_453 = _T_500 ? $signed(dx) : $signed(_GEN_389); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_454 = _T_500 ? $signed(dy) : $signed(_GEN_390); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_455 = _T_500 ? $signed(dz) : $signed(_GEN_391); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_456 = _T_500 ? $signed(dxdx) : $signed(_GEN_392); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_457 = _T_500 ? $signed(dydy) : $signed(_GEN_393); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_458 = _T_500 ? $signed(dzdz) : $signed(_GEN_394); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_459 = _T_500 ? $signed(distance_Reg) : $signed(_GEN_395); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_460 = _T_500 ? $signed(ux) : $signed(_GEN_396); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_461 = _T_500 ? $signed(uy) : $signed(_GEN_397); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_462 = _T_500 ? $signed(uz) : $signed(_GEN_398); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_463 = _T_500 ? $signed(vx) : $signed(_GEN_399); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_464 = _T_500 ? $signed(vy) : $signed(_GEN_400); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_465 = _T_500 ? $signed(vz) : $signed(_GEN_401); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_466 = _T_500 ? $signed(wx) : $signed(_GEN_402); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_467 = _T_500 ? $signed(wy) : $signed(_GEN_403); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_468 = _T_500 ? $signed(wz) : $signed(_GEN_404); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_469 = _T_500 ? $signed(uxux) : $signed(_GEN_405); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_470 = _T_500 ? $signed(uyuy) : $signed(_GEN_406); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_471 = _T_500 ? $signed(uzuz) : $signed(_GEN_407); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_472 = _T_500 ? $signed(uxvx) : $signed(_GEN_408); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_473 = _T_500 ? $signed(uyvy) : $signed(_GEN_409); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_474 = _T_500 ? $signed(uzvz) : $signed(_GEN_410); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_475 = _T_500 ? $signed(vxvx) : $signed(_GEN_411); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_476 = _T_500 ? $signed(vyvy) : $signed(_GEN_412); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_477 = _T_500 ? $signed(vzvz) : $signed(_GEN_413); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_478 = _T_500 ? $signed(uxwx) : $signed(_GEN_414); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_479 = _T_500 ? $signed(uywy) : $signed(_GEN_415); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_480 = _T_500 ? $signed(uzwz) : $signed(_GEN_416); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_481 = _T_500 ? $signed(vxwx) : $signed(_GEN_417); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_482 = _T_500 ? $signed(vywy) : $signed(_GEN_418); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_483 = _T_500 ? $signed(vzwz) : $signed(_GEN_419); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_484 = _T_500 ? $signed(a) : $signed(_GEN_420); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_485 = _T_500 ? $signed(b) : $signed(_GEN_421); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_486 = _T_500 ? $signed(c) : $signed(_GEN_422); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_487 = _T_500 ? $signed(d) : $signed(_GEN_423); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_488 = _T_500 ? $signed(e) : $signed(_GEN_424); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_489 = _T_500 ? $signed(a_ex) : $signed(_GEN_425); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_490 = _T_500 ? $signed(b_ex) : $signed(_GEN_426); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_491 = _T_500 ? $signed(c_ex) : $signed(_GEN_427); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_492 = _T_500 ? $signed(d_ex) : $signed(_GEN_428); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_493 = _T_500 ? $signed(e_ex) : $signed(_GEN_429); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_494 = _T_500 ? $signed(ac) : $signed(_GEN_430); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_495 = _T_500 ? $signed(bb) : $signed(_GEN_431); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_496 = _T_500 ? $signed(be) : $signed(_GEN_432); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_497 = _T_500 ? $signed(cd) : $signed(_GEN_433); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_498 = _T_500 ? $signed(ae) : $signed(_GEN_434); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_499 = _T_500 ? $signed(bd) : $signed(_GEN_435); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_500 = _T_500 ? $signed(D_SUB_B) : $signed(_GEN_436); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_501 = _T_500 ? $signed(sn_temp) : $signed(_GEN_437); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_502 = _T_500 ? $signed(sd_temp) : $signed(_GEN_438); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_503 = _T_500 ? $signed(tn_temp) : $signed(_GEN_439); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_504 = _T_500 ? $signed(td) : $signed(_GEN_440); // @[collide_top.scala 455:9:@545.18]
  assign _GEN_505 = _T_500 ? sd_calData : _GEN_441; // @[collide_top.scala 455:9:@545.18]
  assign _GEN_506 = _T_500 ? td_calData : _GEN_442; // @[collide_top.scala 455:9:@545.18]
  assign _GEN_507 = _T_452 ? {{5'd0}, _T_473} : _GEN_443; // @[collide_top.scala 416:9:@501.16]
  assign _GEN_508 = _T_452 ? {{5'd0}, _T_486} : _GEN_505; // @[collide_top.scala 416:9:@501.16]
  assign _GEN_509 = _T_452 ? {{5'd0}, _T_495} : _GEN_445; // @[collide_top.scala 416:9:@501.16]
  assign _GEN_510 = _T_452 ? {{5'd0}, _T_496} : _GEN_506; // @[collide_top.scala 416:9:@501.16]
  assign _GEN_511 = _T_452 ? 7'h0 : _GEN_444; // @[collide_top.scala 416:9:@501.16]
  assign _GEN_512 = _T_452 ? 7'h0 : _GEN_446; // @[collide_top.scala 416:9:@501.16]
  assign _GEN_513 = _T_452 ? $signed(scux) : $signed(_GEN_447); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_514 = _T_452 ? $signed(tcvx) : $signed(_GEN_448); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_515 = _T_452 ? $signed(scuy) : $signed(_GEN_449); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_516 = _T_452 ? $signed(tcvy) : $signed(_GEN_450); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_517 = _T_452 ? $signed(scuz) : $signed(_GEN_451); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_518 = _T_452 ? $signed(tcvz) : $signed(_GEN_452); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_519 = _T_452 ? $signed(dx) : $signed(_GEN_453); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_520 = _T_452 ? $signed(dy) : $signed(_GEN_454); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_521 = _T_452 ? $signed(dz) : $signed(_GEN_455); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_522 = _T_452 ? $signed(dxdx) : $signed(_GEN_456); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_523 = _T_452 ? $signed(dydy) : $signed(_GEN_457); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_524 = _T_452 ? $signed(dzdz) : $signed(_GEN_458); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_525 = _T_452 ? $signed(distance_Reg) : $signed(_GEN_459); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_526 = _T_452 ? $signed(ux) : $signed(_GEN_460); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_527 = _T_452 ? $signed(uy) : $signed(_GEN_461); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_528 = _T_452 ? $signed(uz) : $signed(_GEN_462); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_529 = _T_452 ? $signed(vx) : $signed(_GEN_463); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_530 = _T_452 ? $signed(vy) : $signed(_GEN_464); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_531 = _T_452 ? $signed(vz) : $signed(_GEN_465); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_532 = _T_452 ? $signed(wx) : $signed(_GEN_466); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_533 = _T_452 ? $signed(wy) : $signed(_GEN_467); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_534 = _T_452 ? $signed(wz) : $signed(_GEN_468); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_535 = _T_452 ? $signed(uxux) : $signed(_GEN_469); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_536 = _T_452 ? $signed(uyuy) : $signed(_GEN_470); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_537 = _T_452 ? $signed(uzuz) : $signed(_GEN_471); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_538 = _T_452 ? $signed(uxvx) : $signed(_GEN_472); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_539 = _T_452 ? $signed(uyvy) : $signed(_GEN_473); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_540 = _T_452 ? $signed(uzvz) : $signed(_GEN_474); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_541 = _T_452 ? $signed(vxvx) : $signed(_GEN_475); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_542 = _T_452 ? $signed(vyvy) : $signed(_GEN_476); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_543 = _T_452 ? $signed(vzvz) : $signed(_GEN_477); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_544 = _T_452 ? $signed(uxwx) : $signed(_GEN_478); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_545 = _T_452 ? $signed(uywy) : $signed(_GEN_479); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_546 = _T_452 ? $signed(uzwz) : $signed(_GEN_480); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_547 = _T_452 ? $signed(vxwx) : $signed(_GEN_481); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_548 = _T_452 ? $signed(vywy) : $signed(_GEN_482); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_549 = _T_452 ? $signed(vzwz) : $signed(_GEN_483); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_550 = _T_452 ? $signed(a) : $signed(_GEN_484); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_551 = _T_452 ? $signed(b) : $signed(_GEN_485); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_552 = _T_452 ? $signed(c) : $signed(_GEN_486); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_553 = _T_452 ? $signed(d) : $signed(_GEN_487); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_554 = _T_452 ? $signed(e) : $signed(_GEN_488); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_555 = _T_452 ? $signed(a_ex) : $signed(_GEN_489); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_556 = _T_452 ? $signed(b_ex) : $signed(_GEN_490); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_557 = _T_452 ? $signed(c_ex) : $signed(_GEN_491); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_558 = _T_452 ? $signed(d_ex) : $signed(_GEN_492); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_559 = _T_452 ? $signed(e_ex) : $signed(_GEN_493); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_560 = _T_452 ? $signed(ac) : $signed(_GEN_494); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_561 = _T_452 ? $signed(bb) : $signed(_GEN_495); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_562 = _T_452 ? $signed(be) : $signed(_GEN_496); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_563 = _T_452 ? $signed(cd) : $signed(_GEN_497); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_564 = _T_452 ? $signed(ae) : $signed(_GEN_498); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_565 = _T_452 ? $signed(bd) : $signed(_GEN_499); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_566 = _T_452 ? $signed(D_SUB_B) : $signed(_GEN_500); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_567 = _T_452 ? $signed(sn_temp) : $signed(_GEN_501); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_568 = _T_452 ? $signed(sd_temp) : $signed(_GEN_502); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_569 = _T_452 ? $signed(tn_temp) : $signed(_GEN_503); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_570 = _T_452 ? $signed(td) : $signed(_GEN_504); // @[collide_top.scala 416:9:@501.16]
  assign _GEN_571 = _T_430 ? $signed(_T_433) : $signed(_GEN_566); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_572 = _T_430 ? $signed(_T_442) : $signed(_GEN_567); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_573 = _T_430 ? $signed(_T_444) : $signed(_GEN_568); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_574 = _T_430 ? $signed(_T_447) : $signed(_GEN_569); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_575 = _T_430 ? $signed(_T_450) : $signed(_GEN_570); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_576 = _T_430 ? sn_calData : _GEN_507; // @[collide_top.scala 388:9:@476.14]
  assign _GEN_577 = _T_430 ? sd_calData : _GEN_508; // @[collide_top.scala 388:9:@476.14]
  assign _GEN_578 = _T_430 ? tn_calData : _GEN_509; // @[collide_top.scala 388:9:@476.14]
  assign _GEN_579 = _T_430 ? td_calData : _GEN_510; // @[collide_top.scala 388:9:@476.14]
  assign _GEN_580 = _T_430 ? {{1'd0}, sc} : _GEN_511; // @[collide_top.scala 388:9:@476.14]
  assign _GEN_581 = _T_430 ? {{1'd0}, tc} : _GEN_512; // @[collide_top.scala 388:9:@476.14]
  assign _GEN_582 = _T_430 ? $signed(scux) : $signed(_GEN_513); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_583 = _T_430 ? $signed(tcvx) : $signed(_GEN_514); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_584 = _T_430 ? $signed(scuy) : $signed(_GEN_515); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_585 = _T_430 ? $signed(tcvy) : $signed(_GEN_516); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_586 = _T_430 ? $signed(scuz) : $signed(_GEN_517); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_587 = _T_430 ? $signed(tcvz) : $signed(_GEN_518); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_588 = _T_430 ? $signed(dx) : $signed(_GEN_519); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_589 = _T_430 ? $signed(dy) : $signed(_GEN_520); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_590 = _T_430 ? $signed(dz) : $signed(_GEN_521); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_591 = _T_430 ? $signed(dxdx) : $signed(_GEN_522); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_592 = _T_430 ? $signed(dydy) : $signed(_GEN_523); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_593 = _T_430 ? $signed(dzdz) : $signed(_GEN_524); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_594 = _T_430 ? $signed(distance_Reg) : $signed(_GEN_525); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_595 = _T_430 ? $signed(ux) : $signed(_GEN_526); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_596 = _T_430 ? $signed(uy) : $signed(_GEN_527); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_597 = _T_430 ? $signed(uz) : $signed(_GEN_528); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_598 = _T_430 ? $signed(vx) : $signed(_GEN_529); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_599 = _T_430 ? $signed(vy) : $signed(_GEN_530); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_600 = _T_430 ? $signed(vz) : $signed(_GEN_531); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_601 = _T_430 ? $signed(wx) : $signed(_GEN_532); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_602 = _T_430 ? $signed(wy) : $signed(_GEN_533); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_603 = _T_430 ? $signed(wz) : $signed(_GEN_534); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_604 = _T_430 ? $signed(uxux) : $signed(_GEN_535); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_605 = _T_430 ? $signed(uyuy) : $signed(_GEN_536); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_606 = _T_430 ? $signed(uzuz) : $signed(_GEN_537); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_607 = _T_430 ? $signed(uxvx) : $signed(_GEN_538); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_608 = _T_430 ? $signed(uyvy) : $signed(_GEN_539); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_609 = _T_430 ? $signed(uzvz) : $signed(_GEN_540); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_610 = _T_430 ? $signed(vxvx) : $signed(_GEN_541); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_611 = _T_430 ? $signed(vyvy) : $signed(_GEN_542); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_612 = _T_430 ? $signed(vzvz) : $signed(_GEN_543); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_613 = _T_430 ? $signed(uxwx) : $signed(_GEN_544); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_614 = _T_430 ? $signed(uywy) : $signed(_GEN_545); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_615 = _T_430 ? $signed(uzwz) : $signed(_GEN_546); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_616 = _T_430 ? $signed(vxwx) : $signed(_GEN_547); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_617 = _T_430 ? $signed(vywy) : $signed(_GEN_548); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_618 = _T_430 ? $signed(vzwz) : $signed(_GEN_549); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_619 = _T_430 ? $signed(a) : $signed(_GEN_550); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_620 = _T_430 ? $signed(b) : $signed(_GEN_551); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_621 = _T_430 ? $signed(c) : $signed(_GEN_552); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_622 = _T_430 ? $signed(d) : $signed(_GEN_553); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_623 = _T_430 ? $signed(e) : $signed(_GEN_554); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_624 = _T_430 ? $signed(a_ex) : $signed(_GEN_555); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_625 = _T_430 ? $signed(b_ex) : $signed(_GEN_556); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_626 = _T_430 ? $signed(c_ex) : $signed(_GEN_557); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_627 = _T_430 ? $signed(d_ex) : $signed(_GEN_558); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_628 = _T_430 ? $signed(e_ex) : $signed(_GEN_559); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_629 = _T_430 ? $signed(ac) : $signed(_GEN_560); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_630 = _T_430 ? $signed(bb) : $signed(_GEN_561); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_631 = _T_430 ? $signed(be) : $signed(_GEN_562); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_632 = _T_430 ? $signed(cd) : $signed(_GEN_563); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_633 = _T_430 ? $signed(ae) : $signed(_GEN_564); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_634 = _T_430 ? $signed(bd) : $signed(_GEN_565); // @[collide_top.scala 388:9:@476.14]
  assign _GEN_635 = _T_382 ? $signed(_T_383) : $signed(_GEN_629); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_636 = _T_382 ? $signed(_T_384) : $signed(_GEN_630); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_637 = _T_382 ? $signed(_T_385) : $signed(_GEN_631); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_638 = _T_382 ? $signed(_T_386) : $signed(_GEN_632); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_639 = _T_382 ? $signed(_T_387) : $signed(_GEN_633); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_640 = _T_382 ? $signed(_T_388) : $signed(_GEN_634); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_641 = _T_382 ? $signed(_T_396) : $signed(_GEN_624); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_642 = _T_382 ? $signed(_T_404) : $signed(_GEN_625); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_643 = _T_382 ? $signed(_T_412) : $signed(_GEN_626); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_644 = _T_382 ? $signed(_T_420) : $signed(_GEN_627); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_645 = _T_382 ? $signed(_T_428) : $signed(_GEN_628); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_646 = _T_382 ? $signed(D_SUB_B) : $signed(_GEN_571); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_647 = _T_382 ? $signed(sn_temp) : $signed(_GEN_572); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_648 = _T_382 ? $signed(sd_temp) : $signed(_GEN_573); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_649 = _T_382 ? $signed(tn_temp) : $signed(_GEN_574); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_650 = _T_382 ? $signed(td) : $signed(_GEN_575); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_651 = _T_382 ? sn_calData : _GEN_576; // @[collide_top.scala 373:9:@425.12]
  assign _GEN_652 = _T_382 ? sd_calData : _GEN_577; // @[collide_top.scala 373:9:@425.12]
  assign _GEN_653 = _T_382 ? tn_calData : _GEN_578; // @[collide_top.scala 373:9:@425.12]
  assign _GEN_654 = _T_382 ? td_calData : _GEN_579; // @[collide_top.scala 373:9:@425.12]
  assign _GEN_655 = _T_382 ? {{1'd0}, sc} : _GEN_580; // @[collide_top.scala 373:9:@425.12]
  assign _GEN_656 = _T_382 ? {{1'd0}, tc} : _GEN_581; // @[collide_top.scala 373:9:@425.12]
  assign _GEN_657 = _T_382 ? $signed(scux) : $signed(_GEN_582); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_658 = _T_382 ? $signed(tcvx) : $signed(_GEN_583); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_659 = _T_382 ? $signed(scuy) : $signed(_GEN_584); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_660 = _T_382 ? $signed(tcvy) : $signed(_GEN_585); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_661 = _T_382 ? $signed(scuz) : $signed(_GEN_586); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_662 = _T_382 ? $signed(tcvz) : $signed(_GEN_587); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_663 = _T_382 ? $signed(dx) : $signed(_GEN_588); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_664 = _T_382 ? $signed(dy) : $signed(_GEN_589); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_665 = _T_382 ? $signed(dz) : $signed(_GEN_590); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_666 = _T_382 ? $signed(dxdx) : $signed(_GEN_591); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_667 = _T_382 ? $signed(dydy) : $signed(_GEN_592); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_668 = _T_382 ? $signed(dzdz) : $signed(_GEN_593); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_669 = _T_382 ? $signed(distance_Reg) : $signed(_GEN_594); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_670 = _T_382 ? $signed(ux) : $signed(_GEN_595); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_671 = _T_382 ? $signed(uy) : $signed(_GEN_596); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_672 = _T_382 ? $signed(uz) : $signed(_GEN_597); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_673 = _T_382 ? $signed(vx) : $signed(_GEN_598); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_674 = _T_382 ? $signed(vy) : $signed(_GEN_599); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_675 = _T_382 ? $signed(vz) : $signed(_GEN_600); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_676 = _T_382 ? $signed(wx) : $signed(_GEN_601); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_677 = _T_382 ? $signed(wy) : $signed(_GEN_602); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_678 = _T_382 ? $signed(wz) : $signed(_GEN_603); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_679 = _T_382 ? $signed(uxux) : $signed(_GEN_604); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_680 = _T_382 ? $signed(uyuy) : $signed(_GEN_605); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_681 = _T_382 ? $signed(uzuz) : $signed(_GEN_606); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_682 = _T_382 ? $signed(uxvx) : $signed(_GEN_607); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_683 = _T_382 ? $signed(uyvy) : $signed(_GEN_608); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_684 = _T_382 ? $signed(uzvz) : $signed(_GEN_609); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_685 = _T_382 ? $signed(vxvx) : $signed(_GEN_610); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_686 = _T_382 ? $signed(vyvy) : $signed(_GEN_611); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_687 = _T_382 ? $signed(vzvz) : $signed(_GEN_612); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_688 = _T_382 ? $signed(uxwx) : $signed(_GEN_613); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_689 = _T_382 ? $signed(uywy) : $signed(_GEN_614); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_690 = _T_382 ? $signed(uzwz) : $signed(_GEN_615); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_691 = _T_382 ? $signed(vxwx) : $signed(_GEN_616); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_692 = _T_382 ? $signed(vywy) : $signed(_GEN_617); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_693 = _T_382 ? $signed(vzwz) : $signed(_GEN_618); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_694 = _T_382 ? $signed(a) : $signed(_GEN_619); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_695 = _T_382 ? $signed(b) : $signed(_GEN_620); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_696 = _T_382 ? $signed(c) : $signed(_GEN_621); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_697 = _T_382 ? $signed(d) : $signed(_GEN_622); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_698 = _T_382 ? $signed(e) : $signed(_GEN_623); // @[collide_top.scala 373:9:@425.12]
  assign _GEN_699 = _T_350 ? $signed(_T_356) : $signed(_GEN_694); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_700 = _T_350 ? $signed(_T_362) : $signed(_GEN_695); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_701 = _T_350 ? $signed(_T_368) : $signed(_GEN_696); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_702 = _T_350 ? $signed(_T_374) : $signed(_GEN_697); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_703 = _T_350 ? $signed(_T_380) : $signed(_GEN_698); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_704 = _T_350 ? $signed(ac) : $signed(_GEN_635); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_705 = _T_350 ? $signed(bb) : $signed(_GEN_636); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_706 = _T_350 ? $signed(be) : $signed(_GEN_637); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_707 = _T_350 ? $signed(cd) : $signed(_GEN_638); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_708 = _T_350 ? $signed(ae) : $signed(_GEN_639); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_709 = _T_350 ? $signed(bd) : $signed(_GEN_640); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_710 = _T_350 ? $signed(a_ex) : $signed(_GEN_641); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_711 = _T_350 ? $signed(b_ex) : $signed(_GEN_642); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_712 = _T_350 ? $signed(c_ex) : $signed(_GEN_643); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_713 = _T_350 ? $signed(d_ex) : $signed(_GEN_644); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_714 = _T_350 ? $signed(e_ex) : $signed(_GEN_645); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_715 = _T_350 ? $signed(D_SUB_B) : $signed(_GEN_646); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_716 = _T_350 ? $signed(sn_temp) : $signed(_GEN_647); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_717 = _T_350 ? $signed(sd_temp) : $signed(_GEN_648); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_718 = _T_350 ? $signed(tn_temp) : $signed(_GEN_649); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_719 = _T_350 ? $signed(td) : $signed(_GEN_650); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_720 = _T_350 ? sn_calData : _GEN_651; // @[collide_top.scala 364:9:@386.10]
  assign _GEN_721 = _T_350 ? sd_calData : _GEN_652; // @[collide_top.scala 364:9:@386.10]
  assign _GEN_722 = _T_350 ? tn_calData : _GEN_653; // @[collide_top.scala 364:9:@386.10]
  assign _GEN_723 = _T_350 ? td_calData : _GEN_654; // @[collide_top.scala 364:9:@386.10]
  assign _GEN_724 = _T_350 ? {{1'd0}, sc} : _GEN_655; // @[collide_top.scala 364:9:@386.10]
  assign _GEN_725 = _T_350 ? {{1'd0}, tc} : _GEN_656; // @[collide_top.scala 364:9:@386.10]
  assign _GEN_726 = _T_350 ? $signed(scux) : $signed(_GEN_657); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_727 = _T_350 ? $signed(tcvx) : $signed(_GEN_658); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_728 = _T_350 ? $signed(scuy) : $signed(_GEN_659); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_729 = _T_350 ? $signed(tcvy) : $signed(_GEN_660); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_730 = _T_350 ? $signed(scuz) : $signed(_GEN_661); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_731 = _T_350 ? $signed(tcvz) : $signed(_GEN_662); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_732 = _T_350 ? $signed(dx) : $signed(_GEN_663); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_733 = _T_350 ? $signed(dy) : $signed(_GEN_664); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_734 = _T_350 ? $signed(dz) : $signed(_GEN_665); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_735 = _T_350 ? $signed(dxdx) : $signed(_GEN_666); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_736 = _T_350 ? $signed(dydy) : $signed(_GEN_667); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_737 = _T_350 ? $signed(dzdz) : $signed(_GEN_668); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_738 = _T_350 ? $signed(distance_Reg) : $signed(_GEN_669); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_739 = _T_350 ? $signed(ux) : $signed(_GEN_670); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_740 = _T_350 ? $signed(uy) : $signed(_GEN_671); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_741 = _T_350 ? $signed(uz) : $signed(_GEN_672); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_742 = _T_350 ? $signed(vx) : $signed(_GEN_673); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_743 = _T_350 ? $signed(vy) : $signed(_GEN_674); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_744 = _T_350 ? $signed(vz) : $signed(_GEN_675); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_745 = _T_350 ? $signed(wx) : $signed(_GEN_676); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_746 = _T_350 ? $signed(wy) : $signed(_GEN_677); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_747 = _T_350 ? $signed(wz) : $signed(_GEN_678); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_748 = _T_350 ? $signed(uxux) : $signed(_GEN_679); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_749 = _T_350 ? $signed(uyuy) : $signed(_GEN_680); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_750 = _T_350 ? $signed(uzuz) : $signed(_GEN_681); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_751 = _T_350 ? $signed(uxvx) : $signed(_GEN_682); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_752 = _T_350 ? $signed(uyvy) : $signed(_GEN_683); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_753 = _T_350 ? $signed(uzvz) : $signed(_GEN_684); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_754 = _T_350 ? $signed(vxvx) : $signed(_GEN_685); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_755 = _T_350 ? $signed(vyvy) : $signed(_GEN_686); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_756 = _T_350 ? $signed(vzvz) : $signed(_GEN_687); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_757 = _T_350 ? $signed(uxwx) : $signed(_GEN_688); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_758 = _T_350 ? $signed(uywy) : $signed(_GEN_689); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_759 = _T_350 ? $signed(uzwz) : $signed(_GEN_690); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_760 = _T_350 ? $signed(vxwx) : $signed(_GEN_691); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_761 = _T_350 ? $signed(vywy) : $signed(_GEN_692); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_762 = _T_350 ? $signed(vzwz) : $signed(_GEN_693); // @[collide_top.scala 364:9:@386.10]
  assign _GEN_763 = _T_333 ? $signed(_T_334) : $signed(_GEN_748); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_764 = _T_333 ? $signed(_T_335) : $signed(_GEN_749); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_765 = _T_333 ? $signed(_T_336) : $signed(_GEN_750); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_766 = _T_333 ? $signed(_T_337) : $signed(_GEN_751); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_767 = _T_333 ? $signed(_T_338) : $signed(_GEN_752); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_768 = _T_333 ? $signed(_T_339) : $signed(_GEN_753); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_769 = _T_333 ? $signed(_T_340) : $signed(_GEN_754); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_770 = _T_333 ? $signed(_T_341) : $signed(_GEN_755); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_771 = _T_333 ? $signed(_T_342) : $signed(_GEN_756); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_772 = _T_333 ? $signed(_T_343) : $signed(_GEN_757); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_773 = _T_333 ? $signed(_T_344) : $signed(_GEN_758); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_774 = _T_333 ? $signed(_T_345) : $signed(_GEN_759); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_775 = _T_333 ? $signed(_T_346) : $signed(_GEN_760); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_776 = _T_333 ? $signed(_T_347) : $signed(_GEN_761); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_777 = _T_333 ? $signed(_T_348) : $signed(_GEN_762); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_778 = _T_333 ? $signed(a) : $signed(_GEN_699); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_779 = _T_333 ? $signed(b) : $signed(_GEN_700); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_780 = _T_333 ? $signed(c) : $signed(_GEN_701); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_781 = _T_333 ? $signed(d) : $signed(_GEN_702); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_782 = _T_333 ? $signed(e) : $signed(_GEN_703); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_783 = _T_333 ? $signed(ac) : $signed(_GEN_704); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_784 = _T_333 ? $signed(bb) : $signed(_GEN_705); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_785 = _T_333 ? $signed(be) : $signed(_GEN_706); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_786 = _T_333 ? $signed(cd) : $signed(_GEN_707); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_787 = _T_333 ? $signed(ae) : $signed(_GEN_708); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_788 = _T_333 ? $signed(bd) : $signed(_GEN_709); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_789 = _T_333 ? $signed(a_ex) : $signed(_GEN_710); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_790 = _T_333 ? $signed(b_ex) : $signed(_GEN_711); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_791 = _T_333 ? $signed(c_ex) : $signed(_GEN_712); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_792 = _T_333 ? $signed(d_ex) : $signed(_GEN_713); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_793 = _T_333 ? $signed(e_ex) : $signed(_GEN_714); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_794 = _T_333 ? $signed(D_SUB_B) : $signed(_GEN_715); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_795 = _T_333 ? $signed(sn_temp) : $signed(_GEN_716); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_796 = _T_333 ? $signed(sd_temp) : $signed(_GEN_717); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_797 = _T_333 ? $signed(tn_temp) : $signed(_GEN_718); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_798 = _T_333 ? $signed(td) : $signed(_GEN_719); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_799 = _T_333 ? sn_calData : _GEN_720; // @[collide_top.scala 346:9:@352.8]
  assign _GEN_800 = _T_333 ? sd_calData : _GEN_721; // @[collide_top.scala 346:9:@352.8]
  assign _GEN_801 = _T_333 ? tn_calData : _GEN_722; // @[collide_top.scala 346:9:@352.8]
  assign _GEN_802 = _T_333 ? td_calData : _GEN_723; // @[collide_top.scala 346:9:@352.8]
  assign _GEN_803 = _T_333 ? {{1'd0}, sc} : _GEN_724; // @[collide_top.scala 346:9:@352.8]
  assign _GEN_804 = _T_333 ? {{1'd0}, tc} : _GEN_725; // @[collide_top.scala 346:9:@352.8]
  assign _GEN_805 = _T_333 ? $signed(scux) : $signed(_GEN_726); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_806 = _T_333 ? $signed(tcvx) : $signed(_GEN_727); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_807 = _T_333 ? $signed(scuy) : $signed(_GEN_728); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_808 = _T_333 ? $signed(tcvy) : $signed(_GEN_729); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_809 = _T_333 ? $signed(scuz) : $signed(_GEN_730); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_810 = _T_333 ? $signed(tcvz) : $signed(_GEN_731); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_811 = _T_333 ? $signed(dx) : $signed(_GEN_732); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_812 = _T_333 ? $signed(dy) : $signed(_GEN_733); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_813 = _T_333 ? $signed(dz) : $signed(_GEN_734); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_814 = _T_333 ? $signed(dxdx) : $signed(_GEN_735); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_815 = _T_333 ? $signed(dydy) : $signed(_GEN_736); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_816 = _T_333 ? $signed(dzdz) : $signed(_GEN_737); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_817 = _T_333 ? $signed(distance_Reg) : $signed(_GEN_738); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_818 = _T_333 ? $signed(ux) : $signed(_GEN_739); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_819 = _T_333 ? $signed(uy) : $signed(_GEN_740); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_820 = _T_333 ? $signed(uz) : $signed(_GEN_741); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_821 = _T_333 ? $signed(vx) : $signed(_GEN_742); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_822 = _T_333 ? $signed(vy) : $signed(_GEN_743); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_823 = _T_333 ? $signed(vz) : $signed(_GEN_744); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_824 = _T_333 ? $signed(wx) : $signed(_GEN_745); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_825 = _T_333 ? $signed(wy) : $signed(_GEN_746); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_826 = _T_333 ? $signed(wz) : $signed(_GEN_747); // @[collide_top.scala 346:9:@352.8]
  assign _GEN_827 = _T_304 ? $signed(_T_307) : $signed(_GEN_818); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_828 = _T_304 ? $signed(_T_310) : $signed(_GEN_819); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_829 = _T_304 ? $signed(_T_313) : $signed(_GEN_820); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_830 = _T_304 ? $signed(_T_316) : $signed(_GEN_821); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_831 = _T_304 ? $signed(_T_319) : $signed(_GEN_822); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_832 = _T_304 ? $signed(_T_322) : $signed(_GEN_823); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_833 = _T_304 ? $signed(_T_325) : $signed(_GEN_824); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_834 = _T_304 ? $signed(_T_328) : $signed(_GEN_825); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_835 = _T_304 ? $signed(_T_331) : $signed(_GEN_826); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_836 = _T_304 ? $signed(uxux) : $signed(_GEN_763); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_837 = _T_304 ? $signed(uyuy) : $signed(_GEN_764); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_838 = _T_304 ? $signed(uzuz) : $signed(_GEN_765); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_839 = _T_304 ? $signed(uxvx) : $signed(_GEN_766); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_840 = _T_304 ? $signed(uyvy) : $signed(_GEN_767); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_841 = _T_304 ? $signed(uzvz) : $signed(_GEN_768); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_842 = _T_304 ? $signed(vxvx) : $signed(_GEN_769); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_843 = _T_304 ? $signed(vyvy) : $signed(_GEN_770); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_844 = _T_304 ? $signed(vzvz) : $signed(_GEN_771); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_845 = _T_304 ? $signed(uxwx) : $signed(_GEN_772); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_846 = _T_304 ? $signed(uywy) : $signed(_GEN_773); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_847 = _T_304 ? $signed(uzwz) : $signed(_GEN_774); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_848 = _T_304 ? $signed(vxwx) : $signed(_GEN_775); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_849 = _T_304 ? $signed(vywy) : $signed(_GEN_776); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_850 = _T_304 ? $signed(vzwz) : $signed(_GEN_777); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_851 = _T_304 ? $signed(a) : $signed(_GEN_778); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_852 = _T_304 ? $signed(b) : $signed(_GEN_779); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_853 = _T_304 ? $signed(c) : $signed(_GEN_780); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_854 = _T_304 ? $signed(d) : $signed(_GEN_781); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_855 = _T_304 ? $signed(e) : $signed(_GEN_782); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_856 = _T_304 ? $signed(ac) : $signed(_GEN_783); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_857 = _T_304 ? $signed(bb) : $signed(_GEN_784); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_858 = _T_304 ? $signed(be) : $signed(_GEN_785); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_859 = _T_304 ? $signed(cd) : $signed(_GEN_786); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_860 = _T_304 ? $signed(ae) : $signed(_GEN_787); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_861 = _T_304 ? $signed(bd) : $signed(_GEN_788); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_862 = _T_304 ? $signed(a_ex) : $signed(_GEN_789); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_863 = _T_304 ? $signed(b_ex) : $signed(_GEN_790); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_864 = _T_304 ? $signed(c_ex) : $signed(_GEN_791); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_865 = _T_304 ? $signed(d_ex) : $signed(_GEN_792); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_866 = _T_304 ? $signed(e_ex) : $signed(_GEN_793); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_867 = _T_304 ? $signed(D_SUB_B) : $signed(_GEN_794); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_868 = _T_304 ? $signed(sn_temp) : $signed(_GEN_795); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_869 = _T_304 ? $signed(sd_temp) : $signed(_GEN_796); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_870 = _T_304 ? $signed(tn_temp) : $signed(_GEN_797); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_871 = _T_304 ? $signed(td) : $signed(_GEN_798); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_872 = _T_304 ? sn_calData : _GEN_799; // @[collide_top.scala 332:9:@312.6]
  assign _GEN_873 = _T_304 ? sd_calData : _GEN_800; // @[collide_top.scala 332:9:@312.6]
  assign _GEN_874 = _T_304 ? tn_calData : _GEN_801; // @[collide_top.scala 332:9:@312.6]
  assign _GEN_875 = _T_304 ? td_calData : _GEN_802; // @[collide_top.scala 332:9:@312.6]
  assign _GEN_876 = _T_304 ? {{1'd0}, sc} : _GEN_803; // @[collide_top.scala 332:9:@312.6]
  assign _GEN_877 = _T_304 ? {{1'd0}, tc} : _GEN_804; // @[collide_top.scala 332:9:@312.6]
  assign _GEN_878 = _T_304 ? $signed(scux) : $signed(_GEN_805); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_879 = _T_304 ? $signed(tcvx) : $signed(_GEN_806); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_880 = _T_304 ? $signed(scuy) : $signed(_GEN_807); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_881 = _T_304 ? $signed(tcvy) : $signed(_GEN_808); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_882 = _T_304 ? $signed(scuz) : $signed(_GEN_809); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_883 = _T_304 ? $signed(tcvz) : $signed(_GEN_810); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_884 = _T_304 ? $signed(dx) : $signed(_GEN_811); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_885 = _T_304 ? $signed(dy) : $signed(_GEN_812); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_886 = _T_304 ? $signed(dz) : $signed(_GEN_813); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_887 = _T_304 ? $signed(dxdx) : $signed(_GEN_814); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_888 = _T_304 ? $signed(dydy) : $signed(_GEN_815); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_889 = _T_304 ? $signed(dzdz) : $signed(_GEN_816); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_890 = _T_304 ? $signed(distance_Reg) : $signed(_GEN_817); // @[collide_top.scala 332:9:@312.6]
  assign _GEN_936 = reset ? 7'h0 : _GEN_876; // @[collide_top.scala 250:1:@244.4]
  assign _GEN_937 = reset ? 7'h0 : _GEN_877; // @[collide_top.scala 250:1:@244.4]
  assign io_distance = distance_Reg; // @[collide_top.scala 590:13:@790.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ux = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  uy = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  uz = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  vx = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  vy = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  vz = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  wx = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  wy = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wz = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  uxux = _RAND_9[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  uyuy = _RAND_10[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  uzuz = _RAND_11[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  uxvx = _RAND_12[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  uyvy = _RAND_13[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  uzvz = _RAND_14[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  vxvx = _RAND_15[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  vyvy = _RAND_16[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  vzvz = _RAND_17[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  uxwx = _RAND_18[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  uywy = _RAND_19[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  uzwz = _RAND_20[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  vxwx = _RAND_21[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  vywy = _RAND_22[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  vzwz = _RAND_23[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  a = _RAND_24[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  b = _RAND_25[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  c = _RAND_26[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  d = _RAND_27[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  e = _RAND_28[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  a_ex = _RAND_29[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  b_ex = _RAND_30[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  c_ex = _RAND_31[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  d_ex = _RAND_32[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  e_ex = _RAND_33[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{`RANDOM}};
  ac = _RAND_34[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  bb = _RAND_35[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  be = _RAND_36[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  cd = _RAND_37[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  ae = _RAND_38[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  bd = _RAND_39[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  D_SUB_B = _RAND_40[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{`RANDOM}};
  sn_temp = _RAND_41[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{`RANDOM}};
  sd_temp = _RAND_42[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  tn_temp = _RAND_43[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {2{`RANDOM}};
  td = _RAND_44[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sc = _RAND_45[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  tc = _RAND_46[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sn_calData = _RAND_47[40:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sd_calData = _RAND_48[40:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  tn_calData = _RAND_49[40:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {2{`RANDOM}};
  td_calData = _RAND_50[40:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  scux = _RAND_51[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  tcvx = _RAND_52[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  scuy = _RAND_53[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  tcvy = _RAND_54[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  scuz = _RAND_55[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  tcvz = _RAND_56[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dx = _RAND_57[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dy = _RAND_58[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dz = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dxdx = _RAND_60[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dydy = _RAND_61[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dzdz = _RAND_62[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  distance_Reg = _RAND_63[17:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ux <= 9'sh0;
    end else begin
      if (_T_304) begin
        ux <= _T_307;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  ux <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uy <= 9'sh0;
    end else begin
      if (_T_304) begin
        uy <= _T_310;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uy <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uz <= 9'sh0;
    end else begin
      if (_T_304) begin
        uz <= _T_313;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uz <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vx <= 9'sh0;
    end else begin
      if (_T_304) begin
        vx <= _T_316;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vx <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vy <= 9'sh0;
    end else begin
      if (_T_304) begin
        vy <= _T_319;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vy <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vz <= 9'sh0;
    end else begin
      if (_T_304) begin
        vz <= _T_322;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vz <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      wx <= 9'sh0;
    end else begin
      if (_T_304) begin
        wx <= _T_325;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  wx <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      wy <= 9'sh0;
    end else begin
      if (_T_304) begin
        wy <= _T_328;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  wy <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      wz <= 9'sh0;
    end else begin
      if (_T_304) begin
        wz <= _T_331;
      end else begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  wz <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uxux <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uxux <= _T_334;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uxux <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uyuy <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uyuy <= _T_335;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uyuy <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uzuz <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uzuz <= _T_336;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uzuz <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uxvx <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uxvx <= _T_337;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uxvx <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uyvy <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uyvy <= _T_338;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uyvy <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uzvz <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uzvz <= _T_339;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uzvz <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vxvx <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          vxvx <= _T_340;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vxvx <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vyvy <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          vyvy <= _T_341;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vyvy <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vzvz <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          vzvz <= _T_342;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vzvz <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uxwx <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uxwx <= _T_343;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uxwx <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uywy <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uywy <= _T_344;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uywy <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      uzwz <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          uzwz <= _T_345;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  uzwz <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vxwx <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          vxwx <= _T_346;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vxwx <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vywy <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          vywy <= _T_347;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vywy <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      vzwz <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (_T_333) begin
          vzwz <= _T_348;
        end else begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  vzwz <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      a <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (_T_350) begin
            a <= _T_356;
          end else begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  a <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      b <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (_T_350) begin
            b <= _T_362;
          end else begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  b <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      c <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (_T_350) begin
            c <= _T_368;
          end else begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  c <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      d <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (_T_350) begin
            d <= _T_374;
          end else begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  d <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      e <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (_T_350) begin
            e <= _T_380;
          end else begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  e <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      a_ex <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              a_ex <= _T_396;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  a_ex <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      b_ex <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              b_ex <= _T_404;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  b_ex <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      c_ex <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              c_ex <= _T_412;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  c_ex <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      d_ex <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              d_ex <= _T_420;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  d_ex <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      e_ex <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              e_ex <= _T_428;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  e_ex <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      ac <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              ac <= _T_383;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  ac <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      bb <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              bb <= _T_384;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  bb <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      be <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              be <= _T_385;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  be <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cd <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              cd <= _T_386;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  cd <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      ae <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              ae <= _T_387;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  ae <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      bd <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (_T_382) begin
              bd <= _T_388;
            end else begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  bd <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      D_SUB_B <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (_T_430) begin
                D_SUB_B <= _T_433;
              end else begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  D_SUB_B <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      sn_temp <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (_T_430) begin
                if (flag_parallel) begin
                  sn_temp <= 36'sh0;
                end else begin
                  if (Foot1OutofSta) begin
                    sn_temp <= 36'sh0;
                  end else begin
                    if (Foot1OutofEnd) begin
                      sn_temp <= _T_439;
                    end else begin
                      sn_temp <= BE_SUB_CD;
                    end
                  end
                end
              end else begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  sn_temp <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      sd_temp <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (_T_430) begin
                if (flag_parallel) begin
                  sd_temp <= 36'sh64;
                end else begin
                  sd_temp <= AC_SUB_BB;
                end
              end else begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  sd_temp <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      tn_temp <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (_T_430) begin
                if (flag_parallel) begin
                  tn_temp <= e_ex;
                end else begin
                  if (Foot1OutofSta) begin
                    tn_temp <= e_ex;
                  end else begin
                    if (Foot1OutofEnd) begin
                      tn_temp <= E_ADD_B;
                    end else begin
                      tn_temp <= AE_SUB_BD;
                    end
                  end
                end
              end else begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  tn_temp <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      td <= 36'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (_T_430) begin
                if (flag_parallel) begin
                  td <= c_ex;
                end else begin
                  if (Foot1OutofSta) begin
                    td <= c_ex;
                  end else begin
                    if (Foot1OutofEnd) begin
                      td <= c_ex;
                    end else begin
                      td <= AC_SUB_BB;
                    end
                  end
                end
              end else begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  td <= 36'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    sc <= _GEN_936[5:0];
    tc <= _GEN_937[5:0];
    if (reset) begin
      sn_calData <= 41'h0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (_T_452) begin
                  sn_calData <= {{5'd0}, _T_473};
                end else begin
                  if (_T_500) begin
                    if (SC_CMP_S2) begin
                      sn_calData <= sn_calData_move2;
                    end else begin
                      sn_calData <= _T_503;
                    end
                  end else begin
                    if (_T_522) begin
                      if (SC_CMP_S2) begin
                        sn_calData <= sn_calData_move2;
                      end else begin
                        sn_calData <= _T_503;
                      end
                    end else begin
                      if (_T_544) begin
                        if (SC_CMP_S2) begin
                          sn_calData <= sn_calData_move2;
                        end else begin
                          sn_calData <= _T_503;
                        end
                      end else begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  sn_calData <= 41'h0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      sd_calData <= 41'h0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (_T_452) begin
                  sd_calData <= {{5'd0}, _T_486};
                end else begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  sd_calData <= 41'h0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      tn_calData <= 41'h0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (_T_452) begin
                  tn_calData <= {{5'd0}, _T_495};
                end else begin
                  if (_T_500) begin
                    if (TC_CMP_S2) begin
                      tn_calData <= tn_calData_move2;
                    end else begin
                      tn_calData <= _T_513;
                    end
                  end else begin
                    if (_T_522) begin
                      if (TC_CMP_S2) begin
                        tn_calData <= tn_calData_move2;
                      end else begin
                        tn_calData <= _T_513;
                      end
                    end else begin
                      if (_T_544) begin
                        if (TC_CMP_S2) begin
                          tn_calData <= tn_calData_move2;
                        end else begin
                          tn_calData <= _T_513;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      td_calData <= 41'h0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (_T_452) begin
                  td_calData <= {{5'd0}, _T_496};
                end else begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  td_calData <= 41'h0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      scux <= 15'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (_T_566) begin
                          scux <= _T_570;
                        end else begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  scux <= 15'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      tcvx <= 15'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (_T_566) begin
                          tcvx <= _T_574;
                        end else begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  tcvx <= 15'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      scuy <= 15'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (_T_566) begin
                          scuy <= _T_578;
                        end else begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  scuy <= 15'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      tcvy <= 15'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (_T_566) begin
                          tcvy <= _T_582;
                        end else begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  tcvy <= 15'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      scuz <= 15'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (_T_566) begin
                          scuz <= _T_586;
                        end else begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  scuz <= 15'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      tcvz <= 15'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (_T_566) begin
                          tcvz <= _T_590;
                        end else begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  tcvz <= 15'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      dx <= 9'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (_T_592) begin
                            dx <= _T_602;
                          end else begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  dx <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      dy <= 9'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (_T_592) begin
                            dy <= _T_612;
                          end else begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  dy <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      dz <= 9'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (_T_592) begin
                            dz <= _T_622;
                          end else begin
                            if (!(_T_624)) begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  dz <= 9'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      dxdx <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (_T_624) begin
                              dxdx <= _T_625;
                            end else begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  dxdx <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      dydy <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (_T_624) begin
                              dydy <= _T_626;
                            end else begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  dydy <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      dzdz <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (_T_624) begin
                              dzdz <= _T_627;
                            end else begin
                              if (!(_T_629)) begin
                                if (!(_T_637)) begin
                                  dzdz <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      distance_Reg <= 18'sh0;
    end else begin
      if (!(_T_304)) begin
        if (!(_T_333)) begin
          if (!(_T_350)) begin
            if (!(_T_382)) begin
              if (!(_T_430)) begin
                if (!(_T_452)) begin
                  if (!(_T_500)) begin
                    if (!(_T_522)) begin
                      if (!(_T_544)) begin
                        if (!(_T_566)) begin
                          if (!(_T_592)) begin
                            if (!(_T_624)) begin
                              if (_T_629) begin
                                distance_Reg <= _T_635;
                              end else begin
                                if (_T_637) begin
                                  distance_Reg <= _T_635;
                                end else begin
                                  distance_Reg <= 18'sh0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
